// Verilog netlist created by TD v5.0.30786
// Wed Aug 24 13:36:24 2022

`timescale 1ns / 1ps
module ROM_Sin_table  // ROM_Sin_table.v(14)
  (
  addra,
  clka,
  rsta,
  doa
  );

  input [15:0] addra;  // ROM_Sin_table.v(18)
  input clka;  // ROM_Sin_table.v(19)
  input rsta;  // ROM_Sin_table.v(20)
  output [11:0] doa;  // ROM_Sin_table.v(16)

  wire [0:2] addra_piped;
  wire  \inst_doa_mux_b0/B0_0 ;
  wire  \inst_doa_mux_b0/B0_1 ;
  wire  \inst_doa_mux_b0/B0_2 ;
  wire  \inst_doa_mux_b0/B0_3 ;
  wire  \inst_doa_mux_b0/B1_0 ;
  wire  \inst_doa_mux_b0/B1_1 ;
  wire  \inst_doa_mux_b1/B0_0 ;
  wire  \inst_doa_mux_b1/B0_1 ;
  wire  \inst_doa_mux_b1/B0_2 ;
  wire  \inst_doa_mux_b1/B0_3 ;
  wire  \inst_doa_mux_b1/B1_0 ;
  wire  \inst_doa_mux_b1/B1_1 ;
  wire  \inst_doa_mux_b10/B0_0 ;
  wire  \inst_doa_mux_b10/B0_1 ;
  wire  \inst_doa_mux_b10/B0_2 ;
  wire  \inst_doa_mux_b10/B0_3 ;
  wire  \inst_doa_mux_b10/B1_0 ;
  wire  \inst_doa_mux_b10/B1_1 ;
  wire  \inst_doa_mux_b11/B0_0 ;
  wire  \inst_doa_mux_b11/B0_1 ;
  wire  \inst_doa_mux_b11/B0_2 ;
  wire  \inst_doa_mux_b11/B0_3 ;
  wire  \inst_doa_mux_b11/B1_0 ;
  wire  \inst_doa_mux_b11/B1_1 ;
  wire  \inst_doa_mux_b2/B0_0 ;
  wire  \inst_doa_mux_b2/B0_1 ;
  wire  \inst_doa_mux_b2/B0_2 ;
  wire  \inst_doa_mux_b2/B0_3 ;
  wire  \inst_doa_mux_b2/B1_0 ;
  wire  \inst_doa_mux_b2/B1_1 ;
  wire  \inst_doa_mux_b3/B0_0 ;
  wire  \inst_doa_mux_b3/B0_1 ;
  wire  \inst_doa_mux_b3/B0_2 ;
  wire  \inst_doa_mux_b3/B0_3 ;
  wire  \inst_doa_mux_b3/B1_0 ;
  wire  \inst_doa_mux_b3/B1_1 ;
  wire  \inst_doa_mux_b4/B0_0 ;
  wire  \inst_doa_mux_b4/B0_1 ;
  wire  \inst_doa_mux_b4/B0_2 ;
  wire  \inst_doa_mux_b4/B0_3 ;
  wire  \inst_doa_mux_b4/B1_0 ;
  wire  \inst_doa_mux_b4/B1_1 ;
  wire  \inst_doa_mux_b5/B0_0 ;
  wire  \inst_doa_mux_b5/B0_1 ;
  wire  \inst_doa_mux_b5/B0_2 ;
  wire  \inst_doa_mux_b5/B0_3 ;
  wire  \inst_doa_mux_b5/B1_0 ;
  wire  \inst_doa_mux_b5/B1_1 ;
  wire  \inst_doa_mux_b6/B0_0 ;
  wire  \inst_doa_mux_b6/B0_1 ;
  wire  \inst_doa_mux_b6/B0_2 ;
  wire  \inst_doa_mux_b6/B0_3 ;
  wire  \inst_doa_mux_b6/B1_0 ;
  wire  \inst_doa_mux_b6/B1_1 ;
  wire  \inst_doa_mux_b7/B0_0 ;
  wire  \inst_doa_mux_b7/B0_1 ;
  wire  \inst_doa_mux_b7/B0_2 ;
  wire  \inst_doa_mux_b7/B0_3 ;
  wire  \inst_doa_mux_b7/B1_0 ;
  wire  \inst_doa_mux_b7/B1_1 ;
  wire  \inst_doa_mux_b8/B0_0 ;
  wire  \inst_doa_mux_b8/B0_1 ;
  wire  \inst_doa_mux_b8/B0_2 ;
  wire  \inst_doa_mux_b8/B0_3 ;
  wire  \inst_doa_mux_b8/B1_0 ;
  wire  \inst_doa_mux_b8/B1_1 ;
  wire  \inst_doa_mux_b9/B0_0 ;
  wire  \inst_doa_mux_b9/B0_1 ;
  wire  \inst_doa_mux_b9/B0_2 ;
  wire  \inst_doa_mux_b9/B0_3 ;
  wire  \inst_doa_mux_b9/B1_0 ;
  wire  \inst_doa_mux_b9/B1_1 ;
  wire inst_doa_i0_000;
  wire inst_doa_i0_001;
  wire inst_doa_i0_002;
  wire inst_doa_i0_003;
  wire inst_doa_i0_004;
  wire inst_doa_i0_005;
  wire inst_doa_i0_006;
  wire inst_doa_i0_007;
  wire inst_doa_i0_008;
  wire inst_doa_i0_009;
  wire inst_doa_i0_010;
  wire inst_doa_i0_011;
  wire inst_doa_i1_000;
  wire inst_doa_i1_001;
  wire inst_doa_i1_002;
  wire inst_doa_i1_003;
  wire inst_doa_i1_004;
  wire inst_doa_i1_005;
  wire inst_doa_i1_006;
  wire inst_doa_i1_007;
  wire inst_doa_i1_008;
  wire inst_doa_i1_009;
  wire inst_doa_i1_010;
  wire inst_doa_i2_000;
  wire inst_doa_i2_001;
  wire inst_doa_i2_002;
  wire inst_doa_i2_003;
  wire inst_doa_i2_004;
  wire inst_doa_i2_005;
  wire inst_doa_i2_006;
  wire inst_doa_i2_007;
  wire inst_doa_i2_008;
  wire inst_doa_i2_009;
  wire inst_doa_i2_010;
  wire inst_doa_i3_000;
  wire inst_doa_i3_001;
  wire inst_doa_i3_002;
  wire inst_doa_i3_003;
  wire inst_doa_i3_004;
  wire inst_doa_i3_005;
  wire inst_doa_i3_006;
  wire inst_doa_i3_007;
  wire inst_doa_i3_008;
  wire inst_doa_i3_009;
  wire inst_doa_i3_010;
  wire inst_doa_i3_011;
  wire inst_doa_i4_000;
  wire inst_doa_i4_001;
  wire inst_doa_i4_002;
  wire inst_doa_i4_003;
  wire inst_doa_i4_004;
  wire inst_doa_i4_005;
  wire inst_doa_i4_006;
  wire inst_doa_i4_007;
  wire inst_doa_i4_008;
  wire inst_doa_i4_009;
  wire inst_doa_i4_010;
  wire inst_doa_i4_011;
  wire inst_doa_i5_000;
  wire inst_doa_i5_001;
  wire inst_doa_i5_002;
  wire inst_doa_i5_003;
  wire inst_doa_i5_004;
  wire inst_doa_i5_005;
  wire inst_doa_i5_006;
  wire inst_doa_i5_007;
  wire inst_doa_i5_008;
  wire inst_doa_i5_009;
  wire inst_doa_i5_010;
  wire inst_doa_i6_000;
  wire inst_doa_i6_001;
  wire inst_doa_i6_002;
  wire inst_doa_i6_003;
  wire inst_doa_i6_004;
  wire inst_doa_i6_005;
  wire inst_doa_i6_006;
  wire inst_doa_i6_007;
  wire inst_doa_i6_008;
  wire inst_doa_i6_009;
  wire inst_doa_i6_010;
  wire inst_doa_i7_000;
  wire inst_doa_i7_001;
  wire inst_doa_i7_002;
  wire inst_doa_i7_003;
  wire inst_doa_i7_004;
  wire inst_doa_i7_005;
  wire inst_doa_i7_006;
  wire inst_doa_i7_007;
  wire inst_doa_i7_008;
  wire inst_doa_i7_009;
  wire inst_doa_i7_010;
  wire inst_doa_i7_011;

  AL_DFF_X addra_pipe_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clka),
    .d(addra[13]),
    .en(1'b1),
    .sr(rsta),
    .ss(1'b0),
    .q(addra_piped[0]));
  AL_DFF_X addra_pipe_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clka),
    .d(addra[14]),
    .en(1'b1),
    .sr(rsta),
    .ss(1'b0),
    .q(addra_piped[1]));
  AL_DFF_X addra_pipe_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clka),
    .d(addra[15]),
    .en(1'b1),
    .sr(rsta),
    .ss(1'b0),
    .q(addra_piped[2]));
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  // address_offset=0;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h7C1F07C1F03E0F83E0F83E0FC1F07C1F07C1F83E0F83E0F83E07C1F07C1F07C0),
    .INIT_01(256'h3E0F83E0FC1F07C1F07C1F83E0F83E0F83F07C1F07C1F07E0F83E0F83E0F81F0),
    .INIT_02(256'h1F07C1F07C0F83E0F83E0F81F07C1F07C1F83E0F83E0F83F07C1F07C1F07E0F8),
    .INIT_03(256'h1F07C0F83E0F83E0FC1F07C1F07C0F83E0F83E0FC1F07C1F07C0F83E0F83E0FC),
    .INIT_04(256'h1F07C1F03E0F83E0F81F07C1F07C0F83E0F83E07C1F07C1F03E0F83E0F81F07C),
    .INIT_05(256'h3E0F83E07C1F07C1F83E0F83E07C1F07C1F83E0F83E07C1F07C1F83E0F83E0FC),
    .INIT_06(256'hF83E0FC1F07C1F83E0F83F07C1F07E0F83E0F81F07C1F03E0F83E07C1F07C1F8),
    .INIT_07(256'hC1F07E0F83E07C1F07C0F83E0FC1F07C0F83E0F81F07C1F03E0F83F07C1F07E0),
    .INIT_08(256'h1F07C0F83E0FC1F07E0F83E07C1F07E0F83E07C1F07E0F83E07C1F07E0F83E07),
    .INIT_09(256'hC1F83E0FC1F07E0F83F07C1F83E0FC1F07C0F83E07C1F03E0F83F07C1F83E0F8),
    .INIT_0A(256'hF81F07C0F83F07C1F83E0FC1F03E0F81F07C0F83F07C1F83E0FC1F07E0F83F07),
    .INIT_0B(256'h7E0F81F07E0F81F07E0F83F07C0F83F07C0F83E07C1F83E07C1F03E0FC1F07E0),
    .INIT_0C(256'h7C0F83F07C0F81F07E0F81F07E0F81F07E0F81F07E0F81F07E0F81F07E0F81F0),
    .INIT_0D(256'hF07E0F81F03E0FC1F83E07C0F83F07E0F81F07E0FC1F03E0FC1F83E07C1F83F0),
    .INIT_0E(256'h0FC1F83F07E0F81F03E07C0F83F07E0FC1F03E07C0F83F07E0FC1F03E07C1F83),
    .INIT_0F(256'hE0FC1F83F07E0FC1F83F07E0FC1F83F07C0F81F03E07C0F81F03E07C0F83F07E),
    .INIT_10(256'hF07E0FC1F81F03E07C0F81F83F07E0FC1F83F03E07C0F81F03E07C0F81F03E07),
    .INIT_11(256'hC1F81F03F07E07C0F81F83F07E07C0F81F83F07E07C0F81F83F07E07C0F81F03),
    .INIT_12(256'h1F83F03E07E0FC0F81F83F03F07E07C0FC1F81F03F07E0FC0F81F83F03E07E0F),
    .INIT_13(256'h83F03F07E07E0FC0FC0F81F81F03F07E07E0FC0FC1F81F83F03E07E07C0FC1F8),
    .INIT_14(256'h81F03F03F03F07E07E07E0FC0FC0F81F81F81F03F03F07E07E07C0FC0F81F81F),
    .INIT_15(256'h1F81F81F81F81F83F03F03F03F03F03E07E07E07E07E0FC0FC0FC0FC1F81F81F),
    .INIT_16(256'hC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0F81F81F8),
    .INIT_17(256'hE07E07E07E03F03F03F03F03F01F81F81F81F81F81F81F80FC0FC0FC0FC0FC0F),
    .INIT_18(256'h03F03F03F81F81F80FC0FC0FE07E07E03F03F03F01F81F81F80FC0FC0FC0FC07),
    .INIT_19(256'hF03F81F80FC0FE07E07F03F01F81FC0FC0FE07E03F03F01F81F80FC0FC07E07E),
    .INIT_1A(256'hF03F81FC0FE07F03F01F80FC0FE07F03F81F80FC0FE07F03F01F81FC0FE07E03),
    .INIT_1B(256'h03F01F80FC07F03F81FC0FE07F01F80FC07E03F01F80FC07E03F01F80FC07E07),
    .INIT_1C(256'hC07E03F80FC07F03F80FC07F03F80FC07F03F80FC07F03F80FC07E03F81FC0FE),
    .INIT_1D(256'h03F80FE03F80FC07F01FC07E03F80FE03F01FC07E03F80FE07F01FC0FE03F81F),
    .INIT_1E(256'hF80FE03F80FE03F80FE03F80FE03F80FE03F80FE03F80FE03F01FC07F01FC07F),
    .INIT_1F(256'hF80FF01FC07F00FE03F80FE03FC07F01FC07F01FC03F80FE03F80FE03F80FE03),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_000000_000 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n66,open_n67,open_n68,open_n69,open_n70,open_n71,open_n72,1'b0,open_n73}),
    .rsta(rsta),
    .doa({open_n88,open_n89,open_n90,open_n91,open_n92,open_n93,open_n94,open_n95,inst_doa_i0_000}));
  // address_offset=0;data_offset=1;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h801FF801FFC00FFC00FFC00FFE007FE007FE003FF003FF003FF801FF801FF800),
    .INIT_01(256'h3FF003FF001FF801FF801FFC00FFC00FFC007FE007FE007FF003FF003FF001FF),
    .INIT_02(256'hE007FE007FF003FF003FF001FF801FF801FFC00FFC00FFC007FE007FE007FF00),
    .INIT_03(256'h1FF800FFC00FFC00FFE007FE007FF003FF003FF001FF801FF800FFC00FFC00FF),
    .INIT_04(256'hE007FE003FF003FF001FF801FF800FFC00FFC007FE007FE003FF003FF001FF80),
    .INIT_05(256'h3FF003FF801FF801FFC00FFC007FE007FE003FF003FF801FF801FFC00FFC00FF),
    .INIT_06(256'h003FF001FF801FFC00FFC007FE007FF003FF001FF801FFC00FFC007FE007FE00),
    .INIT_07(256'hFE007FF003FF801FF800FFC00FFE007FF003FF001FF801FFC00FFC007FE007FF),
    .INIT_08(256'h1FF800FFC00FFE007FF003FF801FF800FFC007FE007FF003FF801FF800FFC007),
    .INIT_09(256'h01FFC00FFE007FF003FF801FFC00FFE007FF003FF801FFC00FFC007FE003FF00),
    .INIT_0A(256'h001FF800FFC007FE003FF001FFC00FFE007FF003FF801FFC00FFE007FF003FF8),
    .INIT_0B(256'h800FFE007FF001FF800FFC007FF003FF800FFC007FE003FF801FFC00FFE007FF),
    .INIT_0C(256'h800FFC007FF001FF800FFE007FF001FF800FFE007FF001FF800FFE007FF001FF),
    .INIT_0D(256'h007FF001FFC00FFE003FF800FFC007FF001FF800FFE003FF001FFC007FE003FF),
    .INIT_0E(256'h0FFE003FF800FFE003FF800FFC007FF001FFC007FF003FF800FFE003FF801FFC),
    .INIT_0F(256'hFF001FFC007FF001FFC007FF001FFC007FF001FFC007FF001FFC007FF003FF80),
    .INIT_10(256'h007FF001FFE003FF800FFE003FF800FFE003FFC007FF001FFC007FF001FFC007),
    .INIT_11(256'hFE001FFC007FF800FFE003FF8007FF001FFC007FF800FFE003FF8007FF001FFC),
    .INIT_12(256'h1FFC003FF800FFF001FFC003FF8007FF001FFE003FF800FFF001FFC003FF800F),
    .INIT_13(256'h03FFC007FF800FFF000FFE001FFC007FF800FFF001FFE003FFC007FF800FFE00),
    .INIT_14(256'h01FFC003FFC007FF8007FF000FFF001FFE001FFC003FF8007FF800FFF001FFE0),
    .INIT_15(256'h1FFE001FFE001FFC003FFC003FFC003FF8007FF8007FF000FFF000FFE001FFE0),
    .INIT_16(256'hFF000FFF000FFF000FFF000FFF000FFF000FFF000FFF000FFF000FFF001FFE00),
    .INIT_17(256'h007FF8007FFC003FFC003FFC001FFE001FFE001FFE001FFF000FFF000FFF000F),
    .INIT_18(256'hFC003FFC001FFE000FFF000FFF8007FFC003FFC001FFE001FFF000FFF000FFF8),
    .INIT_19(256'hFFC001FFF000FFF8007FFC001FFE000FFF0007FFC003FFE001FFF000FFF8007F),
    .INIT_1A(256'hFFC001FFF0007FFC001FFF000FFF8003FFE000FFF0007FFC001FFE000FFF8003),
    .INIT_1B(256'hFC001FFF0007FFC001FFF0007FFE000FFF8003FFE000FFF8003FFE000FFF8007),
    .INIT_1C(256'h007FFC000FFF8003FFF0007FFC000FFF8003FFF0007FFC000FFF8003FFE000FF),
    .INIT_1D(256'hFC000FFFC000FFF8001FFF8003FFF0003FFE0007FFC000FFF8001FFF0003FFE0),
    .INIT_1E(256'hFFF0003FFF0003FFF0003FFF0003FFF0003FFF0003FFF0003FFE0007FFE0007F),
    .INIT_1F(256'hFFF0001FFF8000FFFC000FFFC0007FFE0007FFE0003FFF0003FFF0003FFF0003),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_000000_001 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n124,open_n125,open_n126,open_n127,open_n128,open_n129,open_n130,1'b0,open_n131}),
    .rsta(rsta),
    .doa({open_n146,open_n147,open_n148,open_n149,open_n150,open_n151,open_n152,open_n153,inst_doa_i0_001}));
  // address_offset=0;data_offset=2;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h001FFFFE00000FFFFF00000FFFFF800007FFFFC00003FFFFC00001FFFFE00000),
    .INIT_01(256'hC00003FFFFE00001FFFFE00000FFFFF000007FFFF800007FFFFC00003FFFFE00),
    .INIT_02(256'hFFF800007FFFFC00003FFFFE00001FFFFE00000FFFFF000007FFFF800007FFFF),
    .INIT_03(256'h1FFFFF00000FFFFF000007FFFF800003FFFFC00001FFFFE00000FFFFF00000FF),
    .INIT_04(256'h0007FFFFC00003FFFFE00001FFFFF00000FFFFF800007FFFFC00003FFFFE0000),
    .INIT_05(256'hC00003FFFFE00001FFFFF000007FFFF800003FFFFC00001FFFFE00000FFFFF00),
    .INIT_06(256'hFFC00001FFFFE00000FFFFF800007FFFFC00001FFFFE00000FFFFF800007FFFF),
    .INIT_07(256'hFFFF800003FFFFE00000FFFFF000007FFFFC00001FFFFE00000FFFFF800007FF),
    .INIT_08(256'h1FFFFF00000FFFFF800003FFFFE00000FFFFF800007FFFFC00001FFFFF000007),
    .INIT_09(256'h01FFFFF000007FFFFC00001FFFFF000007FFFFC00001FFFFF000007FFFFC0000),
    .INIT_0A(256'h001FFFFF000007FFFFC00001FFFFF000007FFFFC00001FFFFF000007FFFFC000),
    .INIT_0B(256'h000FFFFF800001FFFFF000007FFFFC00000FFFFF800003FFFFE00000FFFFF800),
    .INIT_0C(256'h000FFFFF800001FFFFF000007FFFFE00000FFFFF800001FFFFF000007FFFFE00),
    .INIT_0D(256'h007FFFFE00000FFFFFC00000FFFFF800001FFFFF000003FFFFE000007FFFFC00),
    .INIT_0E(256'h0FFFFFC00000FFFFFC00000FFFFF800001FFFFF800003FFFFF000003FFFFE000),
    .INIT_0F(256'hFFFFE000007FFFFE000007FFFFE000007FFFFE000007FFFFE000007FFFFC0000),
    .INIT_10(256'hFF800001FFFFFC00000FFFFFC00000FFFFFC000007FFFFE000007FFFFE000007),
    .INIT_11(256'h00001FFFFF800000FFFFFC000007FFFFE000007FFFFF000003FFFFF800001FFF),
    .INIT_12(256'h1FFFFFC00000FFFFFE000003FFFFF800001FFFFFC00000FFFFFE000003FFFFF0),
    .INIT_13(256'hFC000007FFFFF000000FFFFFE000007FFFFF000001FFFFFC000007FFFFF00000),
    .INIT_14(256'h01FFFFFC000007FFFFF800000FFFFFE000001FFFFFC000007FFFFF000001FFFF),
    .INIT_15(256'hE000001FFFFFE000003FFFFFC000003FFFFF8000007FFFFF000000FFFFFE0000),
    .INIT_16(256'hFFFFF000000FFFFFF000000FFFFFF000000FFFFFF000000FFFFFF000001FFFFF),
    .INIT_17(256'h007FFFFF8000003FFFFFC000001FFFFFE000001FFFFFE000000FFFFFF000000F),
    .INIT_18(256'h00003FFFFFE000000FFFFFF0000007FFFFFC000001FFFFFE000000FFFFFF0000),
    .INIT_19(256'h000001FFFFFF0000007FFFFFE000000FFFFFF8000003FFFFFE000000FFFFFF80),
    .INIT_1A(256'h000001FFFFFF8000001FFFFFF0000003FFFFFF0000007FFFFFE000000FFFFFFC),
    .INIT_1B(256'h00001FFFFFF8000001FFFFFF8000000FFFFFFC000000FFFFFFC000000FFFFFF8),
    .INIT_1C(256'h007FFFFFF0000003FFFFFF8000000FFFFFFC0000007FFFFFF0000003FFFFFF00),
    .INIT_1D(256'hFFFFF0000000FFFFFFE0000003FFFFFFC0000007FFFFFF0000001FFFFFFC0000),
    .INIT_1E(256'h0000003FFFFFFC0000003FFFFFFC0000003FFFFFFC0000003FFFFFF80000007F),
    .INIT_1F(256'hFFFFFFE0000000FFFFFFF00000007FFFFFF80000003FFFFFFC0000003FFFFFFC),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_000000_002 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n182,open_n183,open_n184,open_n185,open_n186,open_n187,open_n188,1'b0,open_n189}),
    .rsta(rsta),
    .doa({open_n204,open_n205,open_n206,open_n207,open_n208,open_n209,open_n210,open_n211,inst_doa_i0_002}));
  // address_offset=0;data_offset=3;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h001FFFFFFFFFF0000000000FFFFFFFFFF80000000003FFFFFFFFFE0000000000),
    .INIT_01(256'h000003FFFFFFFFFE0000000000FFFFFFFFFF80000000007FFFFFFFFFC0000000),
    .INIT_02(256'h000000007FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFF80000),
    .INIT_03(256'hE0000000000FFFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF00),
    .INIT_04(256'hFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFF),
    .INIT_05(256'hFFFFFC0000000001FFFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFF),
    .INIT_06(256'hFFFFFFFE0000000000FFFFFFFFFF80000000001FFFFFFFFFF00000000007FFFF),
    .INIT_07(256'hFFFFFFFFFC0000000000FFFFFFFFFF80000000001FFFFFFFFFF00000000007FF),
    .INIT_08(256'h1FFFFFFFFFF00000000003FFFFFFFFFF00000000007FFFFFFFFFE00000000007),
    .INIT_09(256'h01FFFFFFFFFF80000000001FFFFFFFFFF80000000001FFFFFFFFFF8000000000),
    .INIT_0A(256'h001FFFFFFFFFF80000000001FFFFFFFFFF80000000001FFFFFFFFFF800000000),
    .INIT_0B(256'h000FFFFFFFFFFE00000000007FFFFFFFFFF00000000003FFFFFFFFFF00000000),
    .INIT_0C(256'h000FFFFFFFFFFE00000000007FFFFFFFFFF00000000001FFFFFFFFFF80000000),
    .INIT_0D(256'h007FFFFFFFFFF00000000000FFFFFFFFFFE00000000003FFFFFFFFFF80000000),
    .INIT_0E(256'h0FFFFFFFFFFF00000000000FFFFFFFFFFE00000000003FFFFFFFFFFC00000000),
    .INIT_0F(256'hFFFFFFFFFF800000000007FFFFFFFFFF800000000007FFFFFFFFFF8000000000),
    .INIT_10(256'hFFFFFFFE00000000000FFFFFFFFFFF000000000007FFFFFFFFFF800000000007),
    .INIT_11(256'hFFFFE00000000000FFFFFFFFFFF800000000007FFFFFFFFFFC00000000001FFF),
    .INIT_12(256'hE00000000000FFFFFFFFFFFC00000000001FFFFFFFFFFF000000000003FFFFFF),
    .INIT_13(256'h00000007FFFFFFFFFFF000000000007FFFFFFFFFFE000000000007FFFFFFFFFF),
    .INIT_14(256'h01FFFFFFFFFFF800000000000FFFFFFFFFFFE000000000007FFFFFFFFFFE0000),
    .INIT_15(256'hFFFFFFE000000000003FFFFFFFFFFFC000000000007FFFFFFFFFFF0000000000),
    .INIT_16(256'h00000000000FFFFFFFFFFFF000000000000FFFFFFFFFFFF000000000001FFFFF),
    .INIT_17(256'h007FFFFFFFFFFFC000000000001FFFFFFFFFFFE000000000000FFFFFFFFFFFF0),
    .INIT_18(256'hFFFFC000000000000FFFFFFFFFFFF8000000000001FFFFFFFFFFFF0000000000),
    .INIT_19(256'h000001FFFFFFFFFFFF8000000000000FFFFFFFFFFFFC000000000000FFFFFFFF),
    .INIT_1A(256'hFFFFFE0000000000001FFFFFFFFFFFFC0000000000007FFFFFFFFFFFF0000000),
    .INIT_1B(256'h00001FFFFFFFFFFFFE0000000000000FFFFFFFFFFFFF0000000000000FFFFFFF),
    .INIT_1C(256'hFF80000000000003FFFFFFFFFFFFF00000000000007FFFFFFFFFFFFC00000000),
    .INIT_1D(256'hFFFFFFFFFFFF00000000000003FFFFFFFFFFFFF80000000000001FFFFFFFFFFF),
    .INIT_1E(256'h0000003FFFFFFFFFFFFFC00000000000003FFFFFFFFFFFFFC00000000000007F),
    .INIT_1F(256'h00000000000000FFFFFFFFFFFFFF800000000000003FFFFFFFFFFFFFC0000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_000000_003 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n240,open_n241,open_n242,open_n243,open_n244,open_n245,open_n246,1'b0,open_n247}),
    .rsta(rsta),
    .doa({open_n262,open_n263,open_n264,open_n265,open_n266,open_n267,open_n268,open_n269,inst_doa_i0_003}));
  // address_offset=0;data_offset=4;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFE00000000000000000000FFFFFFFFFFFFFFFFFFFFC00000000000000000000),
    .INIT_01(256'h000003FFFFFFFFFFFFFFFFFFFF000000000000000000007FFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFF800000000000000000001FFFFFFFFFFFFFFFFFFFF800000000000000),
    .INIT_03(256'h00000000000FFFFFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFFC000000000),
    .INIT_05(256'h0000000000000001FFFFFFFFFFFFFFFFFFFFC00000000000000000000FFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFF000000000000000000001FFFFFFFFFFFFFFFFFFFF80000),
    .INIT_07(256'h00000000000000000000FFFFFFFFFFFFFFFFFFFFE000000000000000000007FF),
    .INIT_08(256'h1FFFFFFFFFFFFFFFFFFFFC000000000000000000007FFFFFFFFFFFFFFFFFFFF8),
    .INIT_09(256'hFE000000000000000000001FFFFFFFFFFFFFFFFFFFFE00000000000000000000),
    .INIT_0A(256'h001FFFFFFFFFFFFFFFFFFFFE000000000000000000001FFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'hFFF0000000000000000000007FFFFFFFFFFFFFFFFFFFFC000000000000000000),
    .INIT_0C(256'h000FFFFFFFFFFFFFFFFFFFFF8000000000000000000001FFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFF8000000000000000000000FFFFFFFFFFFFFFFFFFFFFC000000000000000000),
    .INIT_0E(256'h0FFFFFFFFFFFFFFFFFFFFFF0000000000000000000003FFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'h0000000000000000000007FFFFFFFFFFFFFFFFFFFFF800000000000000000000),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFF00000000000000000000007FFFFFFFFFFFFFFFFFFFFF8),
    .INIT_11(256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFF80000000000000000000001FFF),
    .INIT_12(256'hFFFFFFFFFFFF00000000000000000000001FFFFFFFFFFFFFFFFFFFFFFC000000),
    .INIT_13(256'h00000007FFFFFFFFFFFFFFFFFFFFFF800000000000000000000007FFFFFFFFFF),
    .INIT_14(256'hFE00000000000000000000000FFFFFFFFFFFFFFFFFFFFFFF8000000000000000),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFC000000000000000000000007FFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'h00000000000FFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000001FFFFF),
    .INIT_17(256'hFF8000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFF0000000000000),
    .INIT_18(256'hFFFFFFFFFFFFFFFFF0000000000000000000000001FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h000001FFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000FFFFFFFF),
    .INIT_1A(256'h0000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000),
    .INIT_1B(256'hFFFFE00000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFF0000000),
    .INIT_1C(256'hFFFFFFFFFFFFFFFC000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000001FFFFFFFFFFF),
    .INIT_1E(256'h0000003FFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000007F),
    .INIT_1F(256'h00000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_000000_004 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n298,open_n299,open_n300,open_n301,open_n302,open_n303,open_n304,1'b0,open_n305}),
    .rsta(rsta),
    .doa({open_n320,open_n321,open_n322,open_n323,open_n324,open_n325,open_n326,open_n327,inst_doa_i0_004}));
  // address_offset=0;data_offset=5;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000),
    .INIT_01(256'hFFFFFC00000000000000000000000000000000000000007FFFFFFFFFFFFFFFFF),
    .INIT_02(256'h00000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'h00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000),
    .INIT_05(256'hFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000FFFFFFF),
    .INIT_06(256'h000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'h00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800),
    .INIT_08(256'h1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000000000),
    .INIT_0A(256'hFFE000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'h0000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'h000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000),
    .INIT_0E(256'hF00000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'h0000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000),
    .INIT_11(256'hFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000001FFF),
    .INIT_12(256'h00000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'h00000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'h00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000000),
    .INIT_18(256'h000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000),
    .INIT_1D(256'h00000000000000000000000000000000000000000000000000001FFFFFFFFFFF),
    .INIT_1E(256'h0000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80),
    .INIT_1F(256'hFFFFFFFFFFFFFF00000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_000000_005 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n356,open_n357,open_n358,open_n359,open_n360,open_n361,open_n362,1'b0,open_n363}),
    .rsta(rsta),
    .doa({open_n378,open_n379,open_n380,open_n381,open_n382,open_n383,open_n384,open_n385,inst_doa_i0_005}));
  // address_offset=0;data_offset=6;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000),
    .INIT_02(256'h00000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFF00000000000000000000000000000000000000000000000000000),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'h000000000000000000000000000000000000000000000000000000000FFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000),
    .INIT_07(256'h00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hE000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'h000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000),
    .INIT_0C(256'h000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000),
    .INIT_0F(256'h0000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000),
    .INIT_12(256'h00000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFF800000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'h0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFFF00000000000000000000000000000000000000000000000000000),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'h000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFE0000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'h0000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000),
    .INIT_1E(256'h0000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_000000_006 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n414,open_n415,open_n416,open_n417,open_n418,open_n419,open_n420,1'b0,open_n421}),
    .rsta(rsta),
    .doa({open_n436,open_n437,open_n438,open_n439,open_n440,open_n441,open_n442,open_n443,inst_doa_i0_006}));
  // address_offset=0;data_offset=7;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'h000000000000000000000000000000000000000000000000000000000FFFFFFF),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'h000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'hFFF0000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'h0000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'h0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'h0000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'hFFFFFFC000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_000000_007 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n472,open_n473,open_n474,open_n475,open_n476,open_n477,open_n478,1'b0,open_n479}),
    .rsta(rsta),
    .doa({open_n494,open_n495,open_n496,open_n497,open_n498,open_n499,open_n500,open_n501,inst_doa_i0_007}));
  // address_offset=0;data_offset=8;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'h000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'h0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_000000_008 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n530,open_n531,open_n532,open_n533,open_n534,open_n535,open_n536,1'b0,open_n537}),
    .rsta(rsta),
    .doa({open_n552,open_n553,open_n554,open_n555,open_n556,open_n557,open_n558,open_n559,inst_doa_i0_008}));
  // address_offset=0;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'h0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_000000_009 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n588,open_n589,open_n590,open_n591,open_n592,open_n593,open_n594,1'b0,open_n595}),
    .rsta(rsta),
    .doa({open_n610,open_n611,open_n612,open_n613,open_n614,open_n615,open_n616,open_n617,inst_doa_i0_009}));
  // address_offset=0;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_000000_010 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n646,open_n647,open_n648,open_n649,open_n650,open_n651,open_n652,1'b0,open_n653}),
    .rsta(rsta),
    .doa({open_n668,open_n669,open_n670,open_n671,open_n672,open_n673,open_n674,open_n675,inst_doa_i0_010}));
  // address_offset=0;data_offset=11;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_000000_011 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n704,open_n705,open_n706,open_n707,open_n708,open_n709,open_n710,1'b0,open_n711}),
    .rsta(rsta),
    .doa({open_n726,open_n727,open_n728,open_n729,open_n730,open_n731,open_n732,open_n733,inst_doa_i0_011}));
  // address_offset=8192;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h03F807F00FE03FC07F00FE03FC07F00FE03F807F01FE03F80FF01FC07F00FE03),
    .INIT_01(256'h00FE01FE03FC07F80FF01FE03FC07F80FF01FE03FC07F80FE01FC03F807F01FE),
    .INIT_02(256'h1FC03FC03F807F807F00FF00FE01FE03FC03F807F80FF00FE01FE03FC07F807F),
    .INIT_03(256'h07F807F807F807F807F807F807F807F807F807F80FF00FF00FF00FE01FE01FE0),
    .INIT_04(256'h7F807F803FC03FC01FE01FE01FF00FF00FF00FF007F807F807F807F807F807F8),
    .INIT_05(256'h0FF807FC03FE01FF00FF807FC03FE01FF00FF007F807FC03FC01FE01FF00FF00),
    .INIT_06(256'hFF007FC01FF00FF803FE01FF007FC03FE00FF007FC03FE00FF007FC03FE01FF0),
    .INIT_07(256'h1FF803FE00FF803FE00FF801FF007FC01FF007FC01FE00FF803FE00FF803FE00),
    .INIT_08(256'hFE007FC00FF801FF003FE007FC01FF803FE007FC01FF803FE00FFC01FF007FC0),
    .INIT_09(256'h7FE007FE007FE007FC00FFC00FFC01FF801FF003FF007FE007FC00FF801FF003),
    .INIT_0A(256'hF801FF800FFC00FFC007FE007FE007FE007FF003FF003FF003FF003FF003FF00),
    .INIT_0B(256'hFE003FF800FFC007FF003FF800FFC007FE003FF801FFC00FFC007FE003FF003F),
    .INIT_0C(256'h007FF800FFE003FFC007FF001FFC007FF001FFC007FF001FFC007FF001FFC007),
    .INIT_0D(256'h003FFC003FFC003FFC007FF8007FF000FFF001FFE003FFC007FF800FFE001FFC),
    .INIT_0E(256'hFFC001FFE000FFF000FFF8007FF8003FFC003FFC003FFC001FFE001FFE001FFE),
    .INIT_0F(256'hFF0007FFE000FFF8003FFE000FFF8003FFE000FFF8007FFC001FFF000FFF8003),
    .INIT_10(256'h0FFFC000FFFC000FFFC000FFFC001FFF8001FFF0003FFF0007FFE000FFF8001F),
    .INIT_11(256'hFFF0001FFFC0007FFF0003FFF8000FFFC0007FFF0003FFF0001FFF8001FFFC00),
    .INIT_12(256'h3FFFC0003FFFC0003FFFC0003FFFC0003FFF80007FFF0000FFFE0003FFF80007),
    .INIT_13(256'hF80001FFFF00003FFFE0000FFFF80003FFFE0001FFFF00007FFF80007FFFC000),
    .INIT_14(256'hFC00007FFFF00003FFFF80000FFFFC0000FFFFC00007FFFE0000FFFFC0000FFF),
    .INIT_15(256'h3FFFFE00000FFFFF800007FFFF800007FFFF800007FFFF80000FFFFE00001FFF),
    .INIT_16(256'hFFFF800000FFFFFE000007FFFFE000003FFFFF000007FFFFE00000FFFFF80000),
    .INIT_17(256'h0FFFFFFC000001FFFFFF0000007FFFFFC000001FFFFFE000001FFFFFC000003F),
    .INIT_18(256'hFFC0000001FFFFFFF00000007FFFFFF80000007FFFFFF0000001FFFFFF800000),
    .INIT_19(256'hFFE000000007FFFFFFFE00000001FFFFFFFE00000001FFFFFFFC0000000FFFFF),
    .INIT_1A(256'h0FFFFFFFFFF8000000000FFFFFFFFFE000000000FFFFFFFFF800000000FFFFFF),
    .INIT_1B(256'hFFFFFFFF0000000000003FFFFFFFFFFF800000000003FFFFFFFFFFC000000000),
    .INIT_1C(256'hFFFFFFFFFFFFFFFE0000000000000007FFFFFFFFFFFFFC00000000000007FFFF),
    .INIT_1D(256'hE000000000000000000000007FFFFFFFFFFFFFFFFFFFE000000000000000000F),
    .INIT_1E(256'h000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_008192_000 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n762,open_n763,open_n764,open_n765,open_n766,open_n767,open_n768,1'b0,open_n769}),
    .rsta(rsta),
    .doa({open_n784,open_n785,open_n786,open_n787,open_n788,open_n789,open_n790,open_n791,inst_doa_i1_000}));
  // address_offset=8192;data_offset=1;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFC0007FFF0003FFF8000FFFC0007FFF0003FFF8001FFFC000FFFE0007FFF0003),
    .INIT_01(256'h00FFFE0003FFF8000FFFE0003FFF8000FFFE0003FFF8000FFFE0003FFF8001FF),
    .INIT_02(256'hE0003FFFC0007FFF8000FFFF0001FFFC0003FFF8000FFFF0001FFFC0007FFF80),
    .INIT_03(256'hF80007FFF80007FFF80007FFF80007FFF80007FFF0000FFFF0000FFFE0001FFF),
    .INIT_04(256'h80007FFFC0003FFFE0001FFFE0000FFFF0000FFFF80007FFF80007FFF80007FF),
    .INIT_05(256'h0FFFF80003FFFE0000FFFF80003FFFE0000FFFF80007FFFC0001FFFE0000FFFF),
    .INIT_06(256'h00007FFFE0000FFFFC0001FFFF80003FFFF00007FFFC0000FFFF80003FFFE000),
    .INIT_07(256'hE00003FFFF00003FFFF00001FFFF80001FFFF80001FFFF00003FFFF00003FFFF),
    .INIT_08(256'h00007FFFF00001FFFFC00007FFFE00003FFFF80001FFFFC0000FFFFE00007FFF),
    .INIT_09(256'h7FFFF800007FFFF80000FFFFF00001FFFFE00003FFFF800007FFFF00001FFFFC),
    .INIT_0A(256'h0001FFFFF00000FFFFF800007FFFF800007FFFFC00003FFFFC00003FFFFC0000),
    .INIT_0B(256'h00003FFFFF000007FFFFC00000FFFFF800003FFFFE00000FFFFF800003FFFFC0),
    .INIT_0C(256'h007FFFFF000003FFFFF800001FFFFF800001FFFFF800001FFFFF800001FFFFF8),
    .INIT_0D(256'hFFC000003FFFFFC000007FFFFF800000FFFFFE000003FFFFF800000FFFFFE000),
    .INIT_0E(256'hFFFFFE000000FFFFFF0000007FFFFFC000003FFFFFC000001FFFFFE000001FFF),
    .INIT_0F(256'hFFFFF8000000FFFFFFC000000FFFFFFC000000FFFFFF8000001FFFFFF0000003),
    .INIT_10(256'hF0000000FFFFFFF0000000FFFFFFE0000001FFFFFFC0000007FFFFFF0000001F),
    .INIT_11(256'hFFFFFFE00000007FFFFFFC0000000FFFFFFF80000003FFFFFFE0000001FFFFFF),
    .INIT_12(256'h3FFFFFFFC00000003FFFFFFFC00000003FFFFFFF80000000FFFFFFFC00000007),
    .INIT_13(256'hFFFFFE000000003FFFFFFFF000000003FFFFFFFE000000007FFFFFFF80000000),
    .INIT_14(256'h0000007FFFFFFFFC000000000FFFFFFFFF0000000007FFFFFFFF000000000FFF),
    .INIT_15(256'hC0000000000FFFFFFFFFF80000000007FFFFFFFFF8000000000FFFFFFFFFE000),
    .INIT_16(256'h0000000000FFFFFFFFFFF800000000003FFFFFFFFFF80000000000FFFFFFFFFF),
    .INIT_17(256'h0FFFFFFFFFFFFE0000000000007FFFFFFFFFFFE000000000001FFFFFFFFFFFC0),
    .INIT_18(256'h0000000001FFFFFFFFFFFFFF800000000000007FFFFFFFFFFFFE000000000000),
    .INIT_19(256'h000000000007FFFFFFFFFFFFFFFE0000000000000001FFFFFFFFFFFFFFF00000),
    .INIT_1A(256'h0FFFFFFFFFFFFFFFFFFFF0000000000000000000FFFFFFFFFFFFFFFFFF000000),
    .INIT_1B(256'h000000000000000000003FFFFFFFFFFFFFFFFFFFFFFC00000000000000000000),
    .INIT_1C(256'h00000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFF80000),
    .INIT_1D(256'h0000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_008192_001 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n820,open_n821,open_n822,open_n823,open_n824,open_n825,open_n826,1'b0,open_n827}),
    .rsta(rsta),
    .doa({open_n842,open_n843,open_n844,open_n845,open_n846,open_n847,open_n848,open_n849,inst_doa_i1_001}));
  // address_offset=8192;data_offset=2;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h000007FFFFFFC0000000FFFFFFF80000003FFFFFFE0000000FFFFFFF80000003),
    .INIT_01(256'hFF00000003FFFFFFF00000003FFFFFFF00000003FFFFFFF00000003FFFFFFE00),
    .INIT_02(256'hFFFFC00000007FFFFFFF00000001FFFFFFFC0000000FFFFFFFE00000007FFFFF),
    .INIT_03(256'hFFFFF800000007FFFFFFF800000007FFFFFFF80000000FFFFFFFF00000001FFF),
    .INIT_04(256'hFFFF800000003FFFFFFFE00000000FFFFFFFF000000007FFFFFFF800000007FF),
    .INIT_05(256'hF000000003FFFFFFFF000000003FFFFFFFF000000007FFFFFFFE00000000FFFF),
    .INIT_06(256'h00007FFFFFFFF000000001FFFFFFFFC000000007FFFFFFFF000000003FFFFFFF),
    .INIT_07(256'hFFFFFC000000003FFFFFFFFE000000001FFFFFFFFE000000003FFFFFFFFC0000),
    .INIT_08(256'h00007FFFFFFFFE0000000007FFFFFFFFC000000001FFFFFFFFF0000000007FFF),
    .INIT_09(256'h80000000007FFFFFFFFF0000000001FFFFFFFFFC0000000007FFFFFFFFE00000),
    .INIT_0A(256'hFFFE0000000000FFFFFFFFFF80000000007FFFFFFFFFC0000000003FFFFFFFFF),
    .INIT_0B(256'hFFFFC00000000007FFFFFFFFFF00000000003FFFFFFFFFF00000000003FFFFFF),
    .INIT_0C(256'hFF800000000003FFFFFFFFFFE00000000001FFFFFFFFFFE00000000001FFFFFF),
    .INIT_0D(256'h000000003FFFFFFFFFFF800000000000FFFFFFFFFFFC00000000000FFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFF0000000000007FFFFFFFFFFFC000000000001FFFFFFFFFFFE000),
    .INIT_0F(256'h000000000000FFFFFFFFFFFFF0000000000000FFFFFFFFFFFFE0000000000003),
    .INIT_10(256'hFFFFFFFF00000000000000FFFFFFFFFFFFFE00000000000007FFFFFFFFFFFFE0),
    .INIT_11(256'hFFFFFFFFFFFFFF800000000000000FFFFFFFFFFFFFFC00000000000001FFFFFF),
    .INIT_12(256'h3FFFFFFFFFFFFFFFC0000000000000003FFFFFFFFFFFFFFF0000000000000007),
    .INIT_13(256'hFFFFFFFFFFFFFFC00000000000000003FFFFFFFFFFFFFFFF8000000000000000),
    .INIT_14(256'hFFFFFF8000000000000000000FFFFFFFFFFFFFFFFFF800000000000000000FFF),
    .INIT_15(256'h00000000000FFFFFFFFFFFFFFFFFFFF80000000000000000000FFFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFF00000000000000000000003FFFFFFFFFFFFFFFFFFFFF0000000000),
    .INIT_17(256'h0FFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000001FFFFFFFFFFFFF),
    .INIT_18(256'h0000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000),
    .INIT_19(256'h000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000),
    .INIT_1A(256'h0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000),
    .INIT_1C(256'h00000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_008192_002 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n878,open_n879,open_n880,open_n881,open_n882,open_n883,open_n884,1'b0,open_n885}),
    .rsta(rsta),
    .doa({open_n900,open_n901,open_n902,open_n903,open_n904,open_n905,open_n906,open_n907,inst_doa_i1_002}));
  // address_offset=8192;data_offset=3;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFF800000000000000FFFFFFFFFFFFFFC00000000000000FFFFFFFFFFFFFFC),
    .INIT_01(256'hFFFFFFFFFC000000000000003FFFFFFFFFFFFFFC000000000000003FFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFF8000000000000001FFFFFFFFFFFFFFF0000000000000007FFFFF),
    .INIT_03(256'hFFFFFFFFFFFFF80000000000000007FFFFFFFFFFFFFFF0000000000000001FFF),
    .INIT_04(256'hFFFFFFFFFFFFC0000000000000000FFFFFFFFFFFFFFFF80000000000000007FF),
    .INIT_05(256'hFFFFFFFFFC00000000000000003FFFFFFFFFFFFFFFF80000000000000000FFFF),
    .INIT_06(256'hFFFF800000000000000001FFFFFFFFFFFFFFFFF800000000000000003FFFFFFF),
    .INIT_07(256'h000000000000003FFFFFFFFFFFFFFFFFE000000000000000003FFFFFFFFFFFFF),
    .INIT_08(256'h00007FFFFFFFFFFFFFFFFFF8000000000000000001FFFFFFFFFFFFFFFFFF8000),
    .INIT_09(256'hFFFFFFFFFF80000000000000000001FFFFFFFFFFFFFFFFFFF800000000000000),
    .INIT_0A(256'h00000000000000FFFFFFFFFFFFFFFFFFFF800000000000000000003FFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFF8000000000000000000003FFFFFFFFFFFFFFFFFFFFC000000),
    .INIT_0C(256'h00000000000003FFFFFFFFFFFFFFFFFFFFFE0000000000000000000001FFFFFF),
    .INIT_0D(256'hFFFFFFFFC00000000000000000000000FFFFFFFFFFFFFFFFFFFFFFF000000000),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000001FFFFFFFFFFFFFFF),
    .INIT_0F(256'h000000000000FFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000003),
    .INIT_10(256'h0000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000),
    .INIT_11(256'h00000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000),
    .INIT_12(256'hC00000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8),
    .INIT_13(256'h00000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'h0000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000),
    .INIT_15(256'h00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000),
    .INIT_17(256'hF00000000000000000000000000000000000000000000000001FFFFFFFFFFFFF),
    .INIT_18(256'h0000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFF80000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_008192_003 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n936,open_n937,open_n938,open_n939,open_n940,open_n941,open_n942,1'b0,open_n943}),
    .rsta(rsta),
    .doa({open_n958,open_n959,open_n960,open_n961,open_n962,open_n963,open_n964,open_n965,inst_doa_i1_003}));
  // address_offset=8192;data_offset=4;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000),
    .INIT_01(256'h0000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000),
    .INIT_02(256'h0000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000),
    .INIT_03(256'h000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000),
    .INIT_04(256'h00000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800),
    .INIT_05(256'h000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000),
    .INIT_06(256'h0000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000),
    .INIT_07(256'h000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000),
    .INIT_08(256'h00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000),
    .INIT_0A(256'hFFFFFFFFFFFFFF00000000000000000000000000000000000000003FFFFFFFFF),
    .INIT_0B(256'h0000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'h00000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFF),
    .INIT_0F(256'h000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000),
    .INIT_11(256'h00000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000),
    .INIT_13(256'h00000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000),
    .INIT_15(256'h00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000),
    .INIT_18(256'h0000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'hF000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_008192_004 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n994,open_n995,open_n996,open_n997,open_n998,open_n999,open_n1000,1'b0,open_n1001}),
    .rsta(rsta),
    .doa({open_n1016,open_n1017,open_n1018,open_n1019,open_n1020,open_n1021,open_n1022,open_n1023,inst_doa_i1_004}));
  // address_offset=8192;data_offset=5;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000),
    .INIT_04(256'h00000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000000),
    .INIT_08(256'h00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000),
    .INIT_0B(256'h0000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFC00000000000000000000000000000000000000000000000000),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFFFF0000000000000000000000000000000000000000000000000000),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h00000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'h00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'hFFFFFFFFFE000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_008192_005 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n1052,open_n1053,open_n1054,open_n1055,open_n1056,open_n1057,open_n1058,1'b0,open_n1059}),
    .rsta(rsta),
    .doa({open_n1074,open_n1075,open_n1076,open_n1077,open_n1078,open_n1079,open_n1080,open_n1081,inst_doa_i1_005}));
  // address_offset=8192;data_offset=6;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'h0000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'h0000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'hFFFF800000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'h0000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h00000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'hFFFFFFFFFFF00000000000000000000000000000000000000000000000000000),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_008192_006 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n1110,open_n1111,open_n1112,open_n1113,open_n1114,open_n1115,open_n1116,1'b0,open_n1117}),
    .rsta(rsta),
    .doa({open_n1132,open_n1133,open_n1134,open_n1135,open_n1136,open_n1137,open_n1138,open_n1139,inst_doa_i1_006}));
  // address_offset=8192;data_offset=7;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'h0000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'h0000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_008192_007 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n1168,open_n1169,open_n1170,open_n1171,open_n1172,open_n1173,open_n1174,1'b0,open_n1175}),
    .rsta(rsta),
    .doa({open_n1190,open_n1191,open_n1192,open_n1193,open_n1194,open_n1195,open_n1196,open_n1197,inst_doa_i1_007}));
  // address_offset=8192;data_offset=8;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'h0000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_008192_008 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n1226,open_n1227,open_n1228,open_n1229,open_n1230,open_n1231,open_n1232,1'b0,open_n1233}),
    .rsta(rsta),
    .doa({open_n1248,open_n1249,open_n1250,open_n1251,open_n1252,open_n1253,open_n1254,open_n1255,inst_doa_i1_008}));
  // address_offset=8192;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_008192_009 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n1284,open_n1285,open_n1286,open_n1287,open_n1288,open_n1289,open_n1290,1'b0,open_n1291}),
    .rsta(rsta),
    .doa({open_n1306,open_n1307,open_n1308,open_n1309,open_n1310,open_n1311,open_n1312,open_n1313,inst_doa_i1_009}));
  // address_offset=8192;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_008192_010 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n1342,open_n1343,open_n1344,open_n1345,open_n1346,open_n1347,open_n1348,1'b0,open_n1349}),
    .rsta(rsta),
    .doa({open_n1364,open_n1365,open_n1366,open_n1367,open_n1368,open_n1369,open_n1370,open_n1371,inst_doa_i1_010}));
  // address_offset=16384;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000),
    .INIT_02(256'hE000000000000000000FFFFFFFFFFFFFFFFFFFFC00000000000000000000000F),
    .INIT_03(256'hFFFFC00000000000007FFFFFFFFFFFFFC000000000000000FFFFFFFFFFFFFFFF),
    .INIT_04(256'h0000000007FFFFFFFFFF800000000003FFFFFFFFFFF8000000000001FFFFFFFF),
    .INIT_05(256'hFFFFFE000000003FFFFFFFFE000000000FFFFFFFFFE0000000003FFFFFFFFFE0),
    .INIT_06(256'hFFFFE00000007FFFFFFF00000000FFFFFFFF00000000FFFFFFFFC00000000FFF),
    .INIT_07(256'h000003FFFFFF0000001FFFFFFC0000003FFFFFFC0000001FFFFFFF00000007FF),
    .INIT_08(256'hF8000007FFFFF000000FFFFFF0000007FFFFFC000001FFFFFF0000007FFFFFE0),
    .INIT_09(256'h00003FFFFE00000FFFFFC00001FFFFF800000FFFFFC00000FFFFFE000003FFFF),
    .INIT_0A(256'hFFF00000FFFFE00003FFFFC00003FFFFC00003FFFFC00003FFFFE00000FFFFF8),
    .INIT_0B(256'hFFE00007FFFE0000FFFFC00007FFFE00007FFFE00003FFFF80001FFFFC00007F),
    .INIT_0C(256'h0007FFFC0003FFFC0001FFFF0000FFFF80003FFFE0000FFFF80001FFFF00003F),
    .INIT_0D(256'hC0003FFF8000FFFE0001FFFC0003FFF80007FFF80007FFF80007FFF80007FFF8),
    .INIT_0E(256'h007FFF0003FFF0001FFF8001FFFC0007FFE0003FFF8001FFFC0007FFF0001FFF),
    .INIT_0F(256'hF0003FFE000FFFC001FFF8001FFF0003FFF0007FFE0007FFE0007FFE0007FFE0),
    .INIT_10(256'h8003FFE001FFF0007FFC003FFE000FFF8003FFE000FFF8003FFE000FFFC001FF),
    .INIT_11(256'hFFF000FFF000FFF0007FF8007FF8007FF8003FFC003FFE001FFE000FFF0007FF),
    .INIT_12(256'h7FF000FFE003FFC007FF800FFF001FFE001FFC003FFC007FF8007FF8007FF800),
    .INIT_13(256'hC007FF001FFC007FF001FFC007FF001FFC007FF001FFC007FF800FFE003FFC00),
    .INIT_14(256'hF801FF800FFC007FE007FF003FF800FFC007FE003FF801FFC007FE003FF800FF),
    .INIT_15(256'h01FF801FF801FF801FF801FF801FFC00FFC00FFC00FFC007FE007FE003FF003F),
    .INIT_16(256'h801FF003FE007FC00FFC01FF801FF003FF007FE007FE007FC00FFC00FFC00FFC),
    .INIT_17(256'h07FC01FF007FE00FF803FF007FC00FF803FF007FC00FF801FF003FE007FC00FF),
    .INIT_18(256'h00FF803FE00FF803FE00FF007FC01FF007FC01FF003FE00FF803FE00FF803FF0),
    .INIT_19(256'h1FF00FF807FC01FE00FF807FC01FE00FF807FC01FF00FF803FE01FF007FC01FE),
    .INIT_1A(256'h01FE01FF00FF007F807FC03FC01FE01FF00FF807FC03FE01FF00FF807FC03FE0),
    .INIT_1B(256'h3FC03FC03FC03FC03FC03FC01FE01FE01FE01FF00FF00FF007F807F803FC03FC),
    .INIT_1C(256'h0FF00FF00FE01FE01FE01FE03FC03FC03FC03FC03FC03FC03FC03FC03FC03FC0),
    .INIT_1D(256'hFC03FC07F80FF00FE01FE03FC03F807F80FF00FE01FE01FC03FC03F807F807F0),
    .INIT_1E(256'hFF01FC03F807F00FE03FC07F80FF01FE03FC07F80FF01FE03FC07F80FF00FE01),
    .INIT_1F(256'h80FE01FC07F01FE03F80FF01FC03F80FE01FC07F80FE01FC07F80FE01FC03F80),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_016384_000 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n1400,open_n1401,open_n1402,open_n1403,open_n1404,open_n1405,open_n1406,1'b0,open_n1407}),
    .rsta(rsta),
    .doa({open_n1422,open_n1423,open_n1424,open_n1425,open_n1426,open_n1427,open_n1428,open_n1429,inst_doa_i2_000}));
  // address_offset=16384;data_offset=1;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'h0000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'h1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000),
    .INIT_03(256'h00003FFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000),
    .INIT_04(256'h000000000000000000007FFFFFFFFFFFFFFFFFFFFFF800000000000000000000),
    .INIT_05(256'h000001FFFFFFFFFFFFFFFFFE0000000000000000001FFFFFFFFFFFFFFFFFFFE0),
    .INIT_06(256'h00001FFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFFC00000000000),
    .INIT_07(256'h000000000000FFFFFFFFFFFFFC00000000000003FFFFFFFFFFFFFF0000000000),
    .INIT_08(256'h07FFFFFFFFFFF000000000000FFFFFFFFFFFFC000000000000FFFFFFFFFFFFE0),
    .INIT_09(256'hFFFFFFFFFE00000000003FFFFFFFFFF800000000003FFFFFFFFFFE0000000000),
    .INIT_0A(256'h000FFFFFFFFFE0000000003FFFFFFFFFC0000000003FFFFFFFFFE00000000007),
    .INIT_0B(256'hFFE000000001FFFFFFFFC000000001FFFFFFFFE0000000007FFFFFFFFC000000),
    .INIT_0C(256'h00000003FFFFFFFC00000000FFFFFFFF800000001FFFFFFFF800000000FFFFFF),
    .INIT_0D(256'hC00000007FFFFFFE00000003FFFFFFF800000007FFFFFFF800000007FFFFFFF8),
    .INIT_0E(256'hFFFFFF0000000FFFFFFF80000003FFFFFFE00000007FFFFFFC0000000FFFFFFF),
    .INIT_0F(256'hF0000001FFFFFFC0000007FFFFFF0000000FFFFFFE0000001FFFFFFE0000001F),
    .INIT_10(256'h8000001FFFFFF0000003FFFFFE0000007FFFFFE0000007FFFFFE0000003FFFFF),
    .INIT_11(256'hFFF000000FFFFFF0000007FFFFF8000007FFFFFC000001FFFFFE000000FFFFFF),
    .INIT_12(256'h000FFFFFE000003FFFFF800000FFFFFE000003FFFFFC000007FFFFF8000007FF),
    .INIT_13(256'h3FFFFF000003FFFFF000003FFFFF000003FFFFF000003FFFFF800001FFFFFC00),
    .INIT_14(256'h07FFFF800003FFFFE00000FFFFF800003FFFFE000007FFFFC00001FFFFF80000),
    .INIT_15(256'h00007FFFF800007FFFF800007FFFFC00003FFFFC00003FFFFE00001FFFFF0000),
    .INIT_16(256'h7FFFF00001FFFFC00003FFFF80000FFFFF00001FFFFE00003FFFFC00003FFFFC),
    .INIT_17(256'hFFFC0000FFFFE00007FFFF00003FFFF80000FFFFC00007FFFF00001FFFFC0000),
    .INIT_18(256'hFFFF80001FFFF80001FFFF00003FFFF00003FFFF00001FFFF80001FFFF80000F),
    .INIT_19(256'h000FFFF80003FFFE00007FFFC0001FFFF80003FFFF00007FFFE0000FFFFC0001),
    .INIT_1A(256'hFFFE0000FFFF00007FFFC0003FFFE0000FFFF80003FFFE0000FFFF80003FFFE0),
    .INIT_1B(256'hFFC0003FFFC0003FFFC0003FFFE0001FFFE0000FFFF0000FFFF80007FFFC0003),
    .INIT_1C(256'hFFF0000FFFE0001FFFE0001FFFC0003FFFC0003FFFC0003FFFC0003FFFC0003F),
    .INIT_1D(256'h03FFFC0007FFF0001FFFE0003FFF80007FFF0001FFFE0003FFFC0007FFF8000F),
    .INIT_1E(256'hFF0003FFF8000FFFE0003FFF8000FFFE0003FFF8000FFFE0003FFF8000FFFE00),
    .INIT_1F(256'h8001FFFC000FFFE0007FFF0003FFF8001FFFC0007FFE0003FFF8001FFFC0007F),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_016384_001 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n1458,open_n1459,open_n1460,open_n1461,open_n1462,open_n1463,open_n1464,1'b0,open_n1465}),
    .rsta(rsta),
    .doa({open_n1480,open_n1481,open_n1482,open_n1483,open_n1484,open_n1485,open_n1486,open_n1487,inst_doa_i2_001}));
  // address_offset=16384;data_offset=2;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'h0000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000),
    .INIT_04(256'h00000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'h000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0),
    .INIT_06(256'h00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000),
    .INIT_07(256'h00000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000),
    .INIT_08(256'hFFFFFFFFFFFFF0000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFE0),
    .INIT_09(256'h0000000001FFFFFFFFFFFFFFFFFFFFF80000000000000000000001FFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFE00000000000000000003FFFFFFFFFFFFFFFFFFFE00000000000),
    .INIT_0B(256'hFFE000000000000000003FFFFFFFFFFFFFFFFFE0000000000000000003FFFFFF),
    .INIT_0C(256'h0000000000000003FFFFFFFFFFFFFFFF800000000000000007FFFFFFFFFFFFFF),
    .INIT_0D(256'hC000000000000001FFFFFFFFFFFFFFF80000000000000007FFFFFFFFFFFFFFF8),
    .INIT_0E(256'hFFFFFF000000000000007FFFFFFFFFFFFFE000000000000003FFFFFFFFFFFFFF),
    .INIT_0F(256'h0FFFFFFFFFFFFFC0000000000000FFFFFFFFFFFFFE00000000000001FFFFFFFF),
    .INIT_10(256'h8000000000000FFFFFFFFFFFFE0000000000001FFFFFFFFFFFFE000000000000),
    .INIT_11(256'h000FFFFFFFFFFFF0000000000007FFFFFFFFFFFC000000000001FFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFE000000000007FFFFFFFFFFE000000000003FFFFFFFFFFF800000000),
    .INIT_13(256'hFFFFFF00000000000FFFFFFFFFFF00000000000FFFFFFFFFFF800000000003FF),
    .INIT_14(256'hFFFFFF80000000001FFFFFFFFFF80000000001FFFFFFFFFFC00000000007FFFF),
    .INIT_15(256'hFFFFFFFFF80000000007FFFFFFFFFC0000000003FFFFFFFFFE0000000000FFFF),
    .INIT_16(256'h00000FFFFFFFFFC0000000007FFFFFFFFF0000000001FFFFFFFFFC0000000003),
    .INIT_17(256'hFFFC000000001FFFFFFFFF0000000007FFFFFFFFC000000000FFFFFFFFFC0000),
    .INIT_18(256'h00007FFFFFFFF800000000FFFFFFFFF000000000FFFFFFFFF8000000007FFFFF),
    .INIT_19(256'hFFFFFFF800000001FFFFFFFFC000000007FFFFFFFF000000001FFFFFFFFC0000),
    .INIT_1A(256'hFFFE00000000FFFFFFFFC00000001FFFFFFFF800000001FFFFFFFF800000001F),
    .INIT_1B(256'hFFC00000003FFFFFFFC00000001FFFFFFFE00000000FFFFFFFF800000003FFFF),
    .INIT_1C(256'hFFF00000001FFFFFFFE00000003FFFFFFFC00000003FFFFFFFC00000003FFFFF),
    .INIT_1D(256'hFFFFFC0000000FFFFFFFE00000007FFFFFFF00000001FFFFFFFC00000007FFFF),
    .INIT_1E(256'h00FFFFFFF80000001FFFFFFF80000001FFFFFFF80000001FFFFFFF80000001FF),
    .INIT_1F(256'h80000003FFFFFFE0000000FFFFFFF80000003FFFFFFE00000007FFFFFFC00000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_016384_002 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n1516,open_n1517,open_n1518,open_n1519,open_n1520,open_n1521,open_n1522,1'b0,open_n1523}),
    .rsta(rsta),
    .doa({open_n1538,open_n1539,open_n1540,open_n1541,open_n1542,open_n1543,open_n1544,open_n1545,inst_doa_i2_002}));
  // address_offset=16384;data_offset=3;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'h000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0),
    .INIT_06(256'h00000000000000000000000000000000000000000000000000003FFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000),
    .INIT_08(256'hFFFFFFFFFFFFF00000000000000000000000000000000000000000000000001F),
    .INIT_09(256'h00000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'h0000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000),
    .INIT_0B(256'h001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000),
    .INIT_0D(256'h3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000007),
    .INIT_0E(256'h000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000),
    .INIT_0F(256'h000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000),
    .INIT_10(256'h80000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFE000000000000),
    .INIT_11(256'hFFFFFFFFFFFFFFF0000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'h000000001FFFFFFFFFFFFFFFFFFFFFFE000000000000000000000007FFFFFFFF),
    .INIT_13(256'hFFFFFF0000000000000000000000FFFFFFFFFFFFFFFFFFFFFF80000000000000),
    .INIT_14(256'h0000007FFFFFFFFFFFFFFFFFFFF8000000000000000000003FFFFFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFF800000000000000000003FFFFFFFFFFFFFFFFFFFE00000000000000),
    .INIT_16(256'h000000000000003FFFFFFFFFFFFFFFFFFF00000000000000000003FFFFFFFFFF),
    .INIT_17(256'h0003FFFFFFFFFFFFFFFFFF0000000000000000003FFFFFFFFFFFFFFFFFFC0000),
    .INIT_18(256'hFFFFFFFFFFFFF800000000000000000FFFFFFFFFFFFFFFFFF800000000000000),
    .INIT_19(256'hFFFFFFF800000000000000003FFFFFFFFFFFFFFFFF000000000000000003FFFF),
    .INIT_1A(256'hFFFE00000000000000003FFFFFFFFFFFFFFFF800000000000000007FFFFFFFFF),
    .INIT_1B(256'hFFC0000000000000003FFFFFFFFFFFFFFFE00000000000000007FFFFFFFFFFFF),
    .INIT_1C(256'hFFF0000000000000001FFFFFFFFFFFFFFFC0000000000000003FFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFC000000000000001FFFFFFFFFFFFFFF0000000000000003FFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFF8000000000000007FFFFFFFFFFFFFF8000000000000007FFFFFFFFF),
    .INIT_1F(256'h7FFFFFFFFFFFFFE000000000000007FFFFFFFFFFFFFE000000000000003FFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_016384_003 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n1574,open_n1575,open_n1576,open_n1577,open_n1578,open_n1579,open_n1580,1'b0,open_n1581}),
    .rsta(rsta),
    .doa({open_n1596,open_n1597,open_n1598,open_n1599,open_n1600,open_n1601,open_n1602,open_n1603,inst_doa_i2_003}));
  // address_offset=16384;data_offset=4;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'h000000000000000000000000000000000000000000000000000000000000001F),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000),
    .INIT_08(256'h0000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000),
    .INIT_0B(256'h000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000),
    .INIT_0D(256'h00000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000),
    .INIT_0F(256'h000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'h7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000),
    .INIT_11(256'hFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000),
    .INIT_12(256'h00000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'h000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000),
    .INIT_15(256'hFFFFFFFFF80000000000000000000000000000000000000001FFFFFFFFFFFFFF),
    .INIT_16(256'h0000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'h0000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000),
    .INIT_18(256'h00000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000),
    .INIT_19(256'h00000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000),
    .INIT_1A(256'h0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000),
    .INIT_1B(256'h003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000),
    .INIT_1C(256'h000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000),
    .INIT_1D(256'h000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000),
    .INIT_1E(256'h0000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000),
    .INIT_1F(256'h000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_016384_004 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n1632,open_n1633,open_n1634,open_n1635,open_n1636,open_n1637,open_n1638,1'b0,open_n1639}),
    .rsta(rsta),
    .doa({open_n1654,open_n1655,open_n1656,open_n1657,open_n1658,open_n1659,open_n1660,open_n1661,inst_doa_i2_004}));
  // address_offset=16384;data_offset=5;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'h000000000000000000000000000000000000000000000000000000FFFFFFFFFF),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'h000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000001FFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'h000000000000000000000000000000000000000000000000007FFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000),
    .INIT_15(256'h0000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000),
    .INIT_18(256'h00000000000000000000000000000000000000000000000007FFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000),
    .INIT_1A(256'h00000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000),
    .INIT_1C(256'h00000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_016384_005 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n1690,open_n1691,open_n1692,open_n1693,open_n1694,open_n1695,open_n1696,1'b0,open_n1697}),
    .rsta(rsta),
    .doa({open_n1712,open_n1713,open_n1714,open_n1715,open_n1716,open_n1717,open_n1718,open_n1719,inst_doa_i2_005}));
  // address_offset=16384;data_offset=6;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'h00000000000000000000000000000000000000000000000000001FFFFFFFFFFF),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'h000000000000000000000000000000000000000000000000000000000003FFFF),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'h00000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'h00000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_016384_006 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n1748,open_n1749,open_n1750,open_n1751,open_n1752,open_n1753,open_n1754,1'b0,open_n1755}),
    .rsta(rsta),
    .doa({open_n1770,open_n1771,open_n1772,open_n1773,open_n1774,open_n1775,open_n1776,open_n1777,inst_doa_i2_006}));
  // address_offset=16384;data_offset=7;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'h00000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_016384_007 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n1806,open_n1807,open_n1808,open_n1809,open_n1810,open_n1811,open_n1812,1'b0,open_n1813}),
    .rsta(rsta),
    .doa({open_n1828,open_n1829,open_n1830,open_n1831,open_n1832,open_n1833,open_n1834,open_n1835,inst_doa_i2_007}));
  // address_offset=16384;data_offset=8;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'h0000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_016384_008 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n1864,open_n1865,open_n1866,open_n1867,open_n1868,open_n1869,open_n1870,1'b0,open_n1871}),
    .rsta(rsta),
    .doa({open_n1886,open_n1887,open_n1888,open_n1889,open_n1890,open_n1891,open_n1892,open_n1893,inst_doa_i2_008}));
  // address_offset=16384;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'h000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_016384_009 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n1922,open_n1923,open_n1924,open_n1925,open_n1926,open_n1927,open_n1928,1'b0,open_n1929}),
    .rsta(rsta),
    .doa({open_n1944,open_n1945,open_n1946,open_n1947,open_n1948,open_n1949,open_n1950,open_n1951,inst_doa_i2_009}));
  // address_offset=16384;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_016384_010 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n1980,open_n1981,open_n1982,open_n1983,open_n1984,open_n1985,open_n1986,1'b0,open_n1987}),
    .rsta(rsta),
    .doa({open_n2002,open_n2003,open_n2004,open_n2005,open_n2006,open_n2007,open_n2008,open_n2009,inst_doa_i2_010}));
  // address_offset=24576;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h80FE03F80FE03F80FE03F807F01FC07F01FC07F80FE03F80FE01FC07F01FE03F),
    .INIT_01(256'hFC07F01FC07F01F80FE03F80FE03F80FE03F80FE03F80FE03F80FE03F80FE03F),
    .INIT_02(256'hF03F80FE07F01FC0FE03F80FC07F01F80FE03F80FC07F01FC07E03F80FE03F81),
    .INIT_03(256'hFE07F03F80FC07E03F81FC07E03F81FC07E03F81FC07E03F81FC07E03F80FC07),
    .INIT_04(256'hC0FC07E03F01F80FC07E03F01F80FC07E03F01FC0FE07F03F81FC07E03F01F80),
    .INIT_05(256'h80FC0FE07F03F01F81FC0FE07E03F03F81FC0FE07E03F01F81FC0FE07F03F81F),
    .INIT_06(256'hFC0FC07E07E03F03F01F81F80FC0FE07E07F03F01F81FC0FC0FE07E03F03F81F),
    .INIT_07(256'hC07E07E07E07E03F03F03F01F81F81F80FC0FC0FE07E07E03F03F03F81F81F80),
    .INIT_08(256'hE07E07E07E07E07E03F03F03F03F03F03F03F01F81F81F81F81F80FC0FC0FC0F),
    .INIT_09(256'h3F03F03E07E07E07E07E07E07E07E07E07E07E07E07E07E07E07E07E07E07E07),
    .INIT_0A(256'hF03F03F07E07E07E07E0FC0FC0FC0FC0F81F81F81F81F81F83F03F03F03F03F0),
    .INIT_0B(256'hF03F03E07E07C0FC0FC1F81F81F03F03F03E07E07E0FC0FC0FC0F81F81F81F03),
    .INIT_0C(256'h3F07E07C0FC0F81F83F03F07E07E0FC0FC1F81F03F03E07E07E0FC0FC1F81F83),
    .INIT_0D(256'hE0FC0F81F83F03E07E0FC1F81F03F07E07C0FC1F81F83F03E07E0FC0F81F83F0),
    .INIT_0E(256'h81F03E07C0FC1F83F03E07C0FC1F83F03E07C0FC1F83F03E07C0FC1F81F03F07),
    .INIT_0F(256'hC0F81F03E07C0F81F03E07C0F81F83F07E0FC1F83F03E07C0F81F03F07E0FC1F),
    .INIT_10(256'hFC1F83E07C0F81F03E07C0F81F03E07C1F83F07E0FC1F83F07E0FC1F83F07E0F),
    .INIT_11(256'h83F07C0F81F07E0FC1F83E07C0F81F07E0FC1F83E07C0F81F03E0FC1F83F07E0),
    .INIT_12(256'h1F83F07C0F83F07E0F81F07E0FC1F03E0FC1F83E07C0F83F07E0F81F03E0FC1F),
    .INIT_13(256'h1F03E0FC1F03E0FC1F03E0FC1F03E0FC1F03E0FC1F03E0FC1F03E07C1F83E07C),
    .INIT_14(256'h0FC1F07E0F81F07C0F83F07C0F83E07C1F83E07C1F83E0FC1F03E0FC1F03E0FC),
    .INIT_15(256'hC1F83E0FC1F07E0F83F07C1F83E07C1F03E0F81F07E0F83F07C1F83E07C1F03E),
    .INIT_16(256'h3E0F83F07C1F83E0F81F07C0F83E07C1F07E0F83F07C1F83E0FC1F07E0F83F07),
    .INIT_17(256'hC0F83E0FC1F07C0F83E0FC1F07C0F83E0FC1F07C0F83E0FC1F07E0F83E07C1F0),
    .INIT_18(256'h0FC1F07C1F83E0F81F07C1F03E0F83E07C1F07E0F83E07C1F07C0F83E0FC1F07),
    .INIT_19(256'h3F07C1F07C0F83E0F81F07C1F03E0F83E0FC1F07C1F83E0F83F07C1F07E0F83E),
    .INIT_1A(256'h7E0F83E0F83F07C1F07C0F83E0F83F07C1F07C0F83E0F83F07C1F07C0F83E0F8),
    .INIT_1B(256'h7C1F03E0F83E0F81F07C1F07C0F83E0F83E07C1F07C1F03E0F83E0F81F07C1F0),
    .INIT_1C(256'h7E0F83E0F83E07C1F07C1F07E0F83E0F83E07C1F07C1F07E0F83E0F83E07C1F0),
    .INIT_1D(256'h3E0FC1F07C1F07C1F83E0F83E0F83F07C1F07C1F03E0F83E0F83E07C1F07C1F0),
    .INIT_1E(256'h1F03E0F83E0F83E0FC1F07C1F07C1F83E0F83E0F83F07C1F07C1F07E0F83E0F8),
    .INIT_1F(256'h07C1F07C1F07C0F83E0F83E0F83F07C1F07C1F07E0F83E0F83E0F81F07C1F07C),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_024576_000 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n2038,open_n2039,open_n2040,open_n2041,open_n2042,open_n2043,open_n2044,1'b0,open_n2045}),
    .rsta(rsta),
    .doa({open_n2060,open_n2061,open_n2062,open_n2063,open_n2064,open_n2065,open_n2066,open_n2067,inst_doa_i3_000}));
  // address_offset=24576;data_offset=1;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h8001FFF8001FFF8001FFF8000FFFC000FFFC0007FFE0007FFE0003FFF0001FFF),
    .INIT_01(256'hFC000FFFC000FFF8001FFF8001FFF8001FFF8001FFF8001FFF8001FFF8001FFF),
    .INIT_02(256'h0FFF8001FFF0003FFE0007FFC000FFF8001FFF8003FFF0003FFE0007FFE0007F),
    .INIT_03(256'hFE000FFF8003FFE0007FFC001FFF8003FFE0007FFC001FFF8003FFE0007FFC00),
    .INIT_04(256'hC003FFE000FFF8003FFE000FFF8003FFE000FFFC001FFF0007FFC001FFF0007F),
    .INIT_05(256'h8003FFE000FFF0007FFC001FFE000FFF8003FFE001FFF0007FFC001FFF0007FF),
    .INIT_06(256'hFC003FFE001FFF000FFF8007FFC001FFE000FFF0007FFC003FFE001FFF0007FF),
    .INIT_07(256'h3FFE001FFE001FFF000FFF0007FF8007FFC003FFE001FFE000FFF0007FF8007F),
    .INIT_08(256'hE001FFE001FFE001FFF000FFF000FFF000FFF0007FF8007FF8007FFC003FFC00),
    .INIT_09(256'h00FFF001FFE001FFE001FFE001FFE001FFE001FFE001FFE001FFE001FFE001FF),
    .INIT_0A(256'h0FFF000FFE001FFE001FFC003FFC003FF8007FF8007FF8007FF000FFF000FFF0),
    .INIT_0B(256'h0FFF001FFE003FFC003FF8007FF000FFF001FFE001FFC003FFC007FF8007FF00),
    .INIT_0C(256'h00FFE003FFC007FF800FFF001FFE003FFC007FF000FFE001FFE003FFC007FF80),
    .INIT_0D(256'hE003FF8007FF001FFE003FF800FFF001FFC003FF8007FF001FFE003FF8007FF0),
    .INIT_0E(256'h7FF001FFC003FF800FFE003FFC007FF001FFC003FF800FFE003FFC007FF000FF),
    .INIT_0F(256'hC007FF001FFC007FF001FFC007FF800FFE003FF800FFE003FF800FFF001FFC00),
    .INIT_10(256'h03FF801FFC007FF001FFC007FF001FFC007FF001FFC007FF001FFC007FF001FF),
    .INIT_11(256'h7FF003FF800FFE003FF801FFC007FF001FFC007FE003FF800FFE003FF800FFE0),
    .INIT_12(256'hFF800FFC007FF001FF800FFE003FF001FFC007FE003FF800FFE007FF001FFC00),
    .INIT_13(256'hFF001FFC00FFE003FF001FFC00FFE003FF001FFC00FFE003FF001FFC007FE003),
    .INIT_14(256'hFFC00FFE007FF003FF800FFC007FE003FF801FFC007FE003FF001FFC00FFE003),
    .INIT_15(256'h3FF801FFC00FFE007FF003FF801FFC00FFE007FF001FF800FFC007FE003FF001),
    .INIT_16(256'h01FF800FFC007FE007FF003FF801FFC00FFE007FF003FF801FFC00FFE007FF00),
    .INIT_17(256'hC007FE003FF003FF801FFC00FFC007FE003FF003FF801FFC00FFE007FE003FF0),
    .INIT_18(256'hFFC00FFC007FE007FF003FF001FF801FFC00FFE007FE003FF003FF801FFC00FF),
    .INIT_19(256'h00FFC00FFC007FE007FF003FF001FF801FFC00FFC007FE007FF003FF001FF801),
    .INIT_1A(256'hFE007FE007FF003FF003FF801FF800FFC00FFC007FE007FF003FF003FF801FF8),
    .INIT_1B(256'h03FF001FF801FF800FFC00FFC007FE007FE003FF003FF001FF801FF800FFC00F),
    .INIT_1C(256'hFE007FE007FE003FF003FF001FF801FF801FFC00FFC00FFE007FE007FE003FF0),
    .INIT_1D(256'h01FFC00FFC00FFC007FE007FE007FF003FF003FF001FF801FF801FFC00FFC00F),
    .INIT_1E(256'hFF001FF801FF801FFC00FFC00FFC007FE007FE007FF003FF003FF001FF801FF8),
    .INIT_1F(256'h003FF003FF003FF801FF801FF800FFC00FFC00FFE007FE007FE007FF003FF003),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_024576_001 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n2096,open_n2097,open_n2098,open_n2099,open_n2100,open_n2101,open_n2102,1'b0,open_n2103}),
    .rsta(rsta),
    .doa({open_n2118,open_n2119,open_n2120,open_n2121,open_n2122,open_n2123,open_n2124,open_n2125,inst_doa_i3_001}));
  // address_offset=24576;data_offset=2;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h7FFFFFF80000007FFFFFF80000003FFFFFFC0000001FFFFFFE0000000FFFFFFF),
    .INIT_01(256'hFC0000003FFFFFF80000007FFFFFF80000007FFFFFF80000007FFFFFF8000000),
    .INIT_02(256'h00007FFFFFF0000001FFFFFFC0000007FFFFFF8000000FFFFFFE0000001FFFFF),
    .INIT_03(256'h01FFFFFF8000001FFFFFFC0000007FFFFFE0000003FFFFFF8000001FFFFFFC00),
    .INIT_04(256'h3FFFFFE0000007FFFFFE0000007FFFFFE0000003FFFFFF0000003FFFFFF00000),
    .INIT_05(256'h7FFFFFE000000FFFFFFC000001FFFFFF8000001FFFFFF0000003FFFFFF000000),
    .INIT_06(256'h03FFFFFE000000FFFFFF8000003FFFFFE000000FFFFFFC000001FFFFFF000000),
    .INIT_07(256'h0001FFFFFE000000FFFFFF0000007FFFFFC000001FFFFFE000000FFFFFF80000),
    .INIT_08(256'hE000001FFFFFE000000FFFFFF000000FFFFFF0000007FFFFF8000003FFFFFC00),
    .INIT_09(256'hFFFFF000001FFFFFE000001FFFFFE000001FFFFFE000001FFFFFE000001FFFFF),
    .INIT_0A(256'h0000FFFFFE000001FFFFFC000003FFFFF8000007FFFFF800000FFFFFF000000F),
    .INIT_0B(256'hFFFF000001FFFFFC000007FFFFF000000FFFFFE000003FFFFFC000007FFFFF00),
    .INIT_0C(256'h00001FFFFFC000007FFFFF000001FFFFFC00000FFFFFE000001FFFFFC000007F),
    .INIT_0D(256'h1FFFFF800000FFFFFE000007FFFFF000003FFFFF800000FFFFFE000007FFFFF0),
    .INIT_0E(256'hFFF000003FFFFF800001FFFFFC00000FFFFFC000007FFFFE000003FFFFF00000),
    .INIT_0F(256'hC00000FFFFFC00000FFFFFC000007FFFFE000007FFFFE000007FFFFF000003FF),
    .INIT_10(256'h00007FFFFC00000FFFFFC00000FFFFFC00000FFFFFC00000FFFFFC00000FFFFF),
    .INIT_11(256'h000FFFFF800001FFFFF800003FFFFF000003FFFFE000007FFFFE000007FFFFE0),
    .INIT_12(256'h007FFFFC00000FFFFF800001FFFFF000003FFFFE000007FFFFE00000FFFFFC00),
    .INIT_13(256'h00FFFFFC00001FFFFF000003FFFFE00000FFFFFC00001FFFFF000003FFFFE000),
    .INIT_14(256'h003FFFFE00000FFFFF800003FFFFE000007FFFFC00001FFFFF000003FFFFE000),
    .INIT_15(256'h0007FFFFC00001FFFFF000007FFFFC00001FFFFF000007FFFFC00001FFFFF000),
    .INIT_16(256'h00007FFFFC00001FFFFF000007FFFFC00001FFFFF000007FFFFC00001FFFFF00),
    .INIT_17(256'hC00001FFFFF000007FFFFC00003FFFFE00000FFFFF800003FFFFE00001FFFFF0),
    .INIT_18(256'hFFC00003FFFFE00000FFFFF000007FFFFC00001FFFFE00000FFFFF800003FFFF),
    .INIT_19(256'hFFFFC00003FFFFE00000FFFFF000007FFFFC00003FFFFE00000FFFFF000007FF),
    .INIT_1A(256'h01FFFFE00000FFFFF000007FFFF800003FFFFC00001FFFFF00000FFFFF800007),
    .INIT_1B(256'h0000FFFFF800007FFFFC00003FFFFE00001FFFFF00000FFFFF800007FFFFC000),
    .INIT_1C(256'hFE00001FFFFE00000FFFFF000007FFFF800003FFFFC00001FFFFE00001FFFFF0),
    .INIT_1D(256'hFFFFC00003FFFFC00001FFFFE00000FFFFF00000FFFFF800007FFFFC00003FFF),
    .INIT_1E(256'h00FFFFF800007FFFFC00003FFFFC00001FFFFE00000FFFFF00000FFFFF800007),
    .INIT_1F(256'h00000FFFFF000007FFFF800007FFFFC00003FFFFE00001FFFFE00000FFFFF000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_024576_002 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n2154,open_n2155,open_n2156,open_n2157,open_n2158,open_n2159,open_n2160,1'b0,open_n2161}),
    .rsta(rsta),
    .doa({open_n2176,open_n2177,open_n2178,open_n2179,open_n2180,open_n2181,open_n2182,open_n2183,inst_doa_i3_002}));
  // address_offset=24576;data_offset=3;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00000007FFFFFFFFFFFFF800000000000003FFFFFFFFFFFFFE00000000000000),
    .INIT_01(256'hFC00000000000007FFFFFFFFFFFFF800000000000007FFFFFFFFFFFFF8000000),
    .INIT_02(256'hFFFFFFFFFFF00000000000003FFFFFFFFFFFFF80000000000001FFFFFFFFFFFF),
    .INIT_03(256'h000000007FFFFFFFFFFFFC0000000000001FFFFFFFFFFFFF80000000000003FF),
    .INIT_04(256'hFFFFFFE0000000000001FFFFFFFFFFFFE0000000000000FFFFFFFFFFFFF00000),
    .INIT_05(256'h0000001FFFFFFFFFFFFC0000000000007FFFFFFFFFFFF0000000000000FFFFFF),
    .INIT_06(256'hFFFFFFFE0000000000007FFFFFFFFFFFE0000000000003FFFFFFFFFFFF000000),
    .INIT_07(256'h0000000001FFFFFFFFFFFF0000000000003FFFFFFFFFFFE0000000000007FFFF),
    .INIT_08(256'h1FFFFFFFFFFFE000000000000FFFFFFFFFFFF0000000000007FFFFFFFFFFFC00),
    .INIT_09(256'hFFFFF000000000001FFFFFFFFFFFE000000000001FFFFFFFFFFFE00000000000),
    .INIT_0A(256'h0000000001FFFFFFFFFFFC000000000007FFFFFFFFFFF800000000000FFFFFFF),
    .INIT_0B(256'h0000FFFFFFFFFFFC00000000000FFFFFFFFFFFE000000000003FFFFFFFFFFF00),
    .INIT_0C(256'hFFFFFFFFFFC00000000000FFFFFFFFFFFC00000000001FFFFFFFFFFFC0000000),
    .INIT_0D(256'hFFFFFF800000000001FFFFFFFFFFF000000000007FFFFFFFFFFE00000000000F),
    .INIT_0E(256'hFFF000000000007FFFFFFFFFFC00000000003FFFFFFFFFFE00000000000FFFFF),
    .INIT_0F(256'hC00000000003FFFFFFFFFFC00000000001FFFFFFFFFFE00000000000FFFFFFFF),
    .INIT_10(256'h0000000003FFFFFFFFFFC00000000003FFFFFFFFFFC00000000003FFFFFFFFFF),
    .INIT_11(256'h000000007FFFFFFFFFF80000000000FFFFFFFFFFE00000000001FFFFFFFFFFE0),
    .INIT_12(256'h00000003FFFFFFFFFF80000000000FFFFFFFFFFE00000000001FFFFFFFFFFC00),
    .INIT_13(256'h00000003FFFFFFFFFF00000000001FFFFFFFFFFC0000000000FFFFFFFFFFE000),
    .INIT_14(256'h00000001FFFFFFFFFF80000000001FFFFFFFFFFC0000000000FFFFFFFFFFE000),
    .INIT_15(256'h000000003FFFFFFFFFF00000000003FFFFFFFFFF00000000003FFFFFFFFFF000),
    .INIT_16(256'h0000000003FFFFFFFFFF00000000003FFFFFFFFFF00000000003FFFFFFFFFF00),
    .INIT_17(256'hC0000000000FFFFFFFFFFC0000000001FFFFFFFFFF80000000001FFFFFFFFFF0),
    .INIT_18(256'hFFC0000000001FFFFFFFFFF00000000003FFFFFFFFFE00000000007FFFFFFFFF),
    .INIT_19(256'hFFFFC0000000001FFFFFFFFFF00000000003FFFFFFFFFE0000000000FFFFFFFF),
    .INIT_1A(256'hFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFFF00000000007FFFFF),
    .INIT_1B(256'hFFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFF),
    .INIT_1C(256'h01FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFFFE0000000000F),
    .INIT_1D(256'h00003FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFFC00000000),
    .INIT_1E(256'h00000007FFFFFFFFFC0000000003FFFFFFFFFE0000000000FFFFFFFFFF800000),
    .INIT_1F(256'h0000000000FFFFFFFFFF80000000003FFFFFFFFFE0000000001FFFFFFFFFF000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_024576_003 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n2212,open_n2213,open_n2214,open_n2215,open_n2216,open_n2217,open_n2218,1'b0,open_n2219}),
    .rsta(rsta),
    .doa({open_n2234,open_n2235,open_n2236,open_n2237,open_n2238,open_n2239,open_n2240,open_n2241,inst_doa_i3_003}));
  // address_offset=24576;data_offset=4;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000),
    .INIT_01(256'hFC0000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFF8000000),
    .INIT_02(256'hFFFFFFFFFFF0000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000007FFFFFFFFFFFFFFF),
    .INIT_04(256'h0000001FFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000FFFFF),
    .INIT_05(256'h00000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000),
    .INIT_06(256'hFFFFFFFE0000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFF000000),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000001FFFFFFFFFFFFFFFFF),
    .INIT_08(256'h0000000000001FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000003FF),
    .INIT_09(256'hFFFFF000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFE00000000000),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFC000000000000000000000007FFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'h0000000000000003FFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000FF),
    .INIT_0C(256'hFFFFFFFFFFC00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFC0000000),
    .INIT_0D(256'h0000007FFFFFFFFFFFFFFFFFFFFFF00000000000000000000001FFFFFFFFFFFF),
    .INIT_0E(256'hFFF00000000000000000000003FFFFFFFFFFFFFFFFFFFFFE0000000000000000),
    .INIT_0F(256'h3FFFFFFFFFFFFFFFFFFFFFC0000000000000000000001FFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'h000000000000000000003FFFFFFFFFFFFFFFFFFFFFC000000000000000000000),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFF8000000000000000000001FFFFFFFFFFFFFFFFFFFFFE0),
    .INIT_12(256'h0000000000000000007FFFFFFFFFFFFFFFFFFFFE0000000000000000000003FF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFF0000000000000000000003FFFFFFFFFFFFFFFFFFFFE000),
    .INIT_14(256'h0000000000000000007FFFFFFFFFFFFFFFFFFFFC000000000000000000001FFF),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFF000000000000000000000FFFFFFFFFFFFFFFFFFFFF000),
    .INIT_16(256'h00000000000000000000FFFFFFFFFFFFFFFFFFFFF000000000000000000000FF),
    .INIT_17(256'h3FFFFFFFFFFFFFFFFFFFFC000000000000000000007FFFFFFFFFFFFFFFFFFFF0),
    .INIT_18(256'hFFC00000000000000000000FFFFFFFFFFFFFFFFFFFFE00000000000000000000),
    .INIT_19(256'h00003FFFFFFFFFFFFFFFFFFFF000000000000000000001FFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFE000000000000000000007FFFFFFFFFFFFFFFFFFFF0000000000000000),
    .INIT_1B(256'h0000000007FFFFFFFFFFFFFFFFFFFE000000000000000000007FFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFE000000000000000000007FFFFFFFFFFFFFFFFFFFE00000000000),
    .INIT_1D(256'h000000000000003FFFFFFFFFFFFFFFFFFFF000000000000000000003FFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFC00000000000000000001FFFFFFFFFFFFFFFFFFFF800000),
    .INIT_1F(256'h000000000000000000007FFFFFFFFFFFFFFFFFFFE00000000000000000000FFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_024576_004 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n2270,open_n2271,open_n2272,open_n2273,open_n2274,open_n2275,open_n2276,1'b0,open_n2277}),
    .rsta(rsta),
    .doa({open_n2292,open_n2293,open_n2294,open_n2295,open_n2296,open_n2297,open_n2298,open_n2299,inst_doa_i3_004}));
  // address_offset=24576;data_offset=5;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00000000000000000000000000000000000000000000000001FFFFFFFFFFFFFF),
    .INIT_01(256'h03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000),
    .INIT_02(256'hFFFFFFFFFFF00000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000),
    .INIT_05(256'h000000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'h00000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'h00000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000),
    .INIT_0B(256'h000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'h00000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000),
    .INIT_0E(256'hFFF000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFF),
    .INIT_0F(256'h00000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000000000000001F),
    .INIT_12(256'h0000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'h000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000FFF),
    .INIT_16(256'h00000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'h0000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0),
    .INIT_18(256'h003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000),
    .INIT_1A(256'hFFFFFFE00000000000000000000000000000000000000000FFFFFFFFFFFFFFFF),
    .INIT_1B(256'h000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'h000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000007FFFFF),
    .INIT_1F(256'h00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_024576_005 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n2328,open_n2329,open_n2330,open_n2331,open_n2332,open_n2333,open_n2334,1'b0,open_n2335}),
    .rsta(rsta),
    .doa({open_n2350,open_n2351,open_n2352,open_n2353,open_n2354,open_n2355,open_n2356,open_n2357,inst_doa_i3_005}));
  // address_offset=24576;data_offset=6;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000),
    .INIT_02(256'h00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000FFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'h00000000000000000000000000000000000000000000000000001FFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'h000000000000000000000000000000000000000000000000000000003FFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000),
    .INIT_0E(256'h000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000),
    .INIT_11(256'h00000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000),
    .INIT_14(256'h0000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'h000000000000000000000000000000000000000000000000000000000000000F),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000),
    .INIT_19(256'h0000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFE000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'h00000000000000000000000000000000000000000000000000001FFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000),
    .INIT_1E(256'h000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_024576_006 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n2386,open_n2387,open_n2388,open_n2389,open_n2390,open_n2391,open_n2392,1'b0,open_n2393}),
    .rsta(rsta),
    .doa({open_n2408,open_n2409,open_n2410,open_n2411,open_n2412,open_n2413,open_n2414,open_n2415,inst_doa_i3_006}));
  // address_offset=24576;data_offset=7;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000007FFFFFF),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'h0000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'h00000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000001FFF),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'h00000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'hFFFFFFE000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'h00000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_024576_007 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n2444,open_n2445,open_n2446,open_n2447,open_n2448,open_n2449,open_n2450,1'b0,open_n2451}),
    .rsta(rsta),
    .doa({open_n2466,open_n2467,open_n2468,open_n2469,open_n2470,open_n2471,open_n2472,open_n2473,inst_doa_i3_007}));
  // address_offset=24576;data_offset=8;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'h000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'h0000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'h0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_024576_008 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n2502,open_n2503,open_n2504,open_n2505,open_n2506,open_n2507,open_n2508,1'b0,open_n2509}),
    .rsta(rsta),
    .doa({open_n2524,open_n2525,open_n2526,open_n2527,open_n2528,open_n2529,open_n2530,open_n2531,inst_doa_i3_008}));
  // address_offset=24576;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'h0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_024576_009 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n2560,open_n2561,open_n2562,open_n2563,open_n2564,open_n2565,open_n2566,1'b0,open_n2567}),
    .rsta(rsta),
    .doa({open_n2582,open_n2583,open_n2584,open_n2585,open_n2586,open_n2587,open_n2588,open_n2589,inst_doa_i3_009}));
  // address_offset=24576;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'h0000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_024576_010 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n2618,open_n2619,open_n2620,open_n2621,open_n2622,open_n2623,open_n2624,1'b0,open_n2625}),
    .rsta(rsta),
    .doa({open_n2640,open_n2641,open_n2642,open_n2643,open_n2644,open_n2645,open_n2646,open_n2647,inst_doa_i3_010}));
  // address_offset=24576;data_offset=11;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_024576_011 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n2676,open_n2677,open_n2678,open_n2679,open_n2680,open_n2681,open_n2682,1'b0,open_n2683}),
    .rsta(rsta),
    .doa({open_n2698,open_n2699,open_n2700,open_n2701,open_n2702,open_n2703,open_n2704,open_n2705,inst_doa_i3_011}));
  // address_offset=32768;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h83E0F83E0FC1F07C1F07C1F03E0F83E0F83E07C1F07C1F07C1F83E0F83E0F83F),
    .INIT_01(256'hC1F07C1F03E0F83E0F83E07C1F07C1F07C0F83E0F83E0F81F07C1F07C1F07E0F),
    .INIT_02(256'hE0F83E0F83F07C1F07C1F07E0F83E0F83E07C1F07C1F07C0F83E0F83E0F81F07),
    .INIT_03(256'hE0F83F07C1F07C1F03E0F83E0F83F07C1F07C1F03E0F83E0F83F07C1F07C1F03),
    .INIT_04(256'hE0F83E0FC1F07C1F07E0F83E0F83F07C1F07C1F83E0F83E0FC1F07C1F07E0F83),
    .INIT_05(256'hC1F07C1F83E0F83E07C1F07C1F83E0F83E07C1F07C1F83E0F83E07C1F07C1F03),
    .INIT_06(256'h07C1F03E0F83E07C1F07C0F83E0F81F07C1F07E0F83E0FC1F07C1F83E0F83E07),
    .INIT_07(256'h3E0F81F07C1F83E0F83F07C1F03E0F83F07C1F07E0F83E0FC1F07C0F83E0F81F),
    .INIT_08(256'hE0F83F07C1F03E0F81F07C1F83E0F81F07C1F83E0F81F07C1F83E0F81F07C1F8),
    .INIT_09(256'h3E07C1F03E0F81F07C0F83E07C1F03E0F83F07C1F83E0FC1F07C0F83E07C1F07),
    .INIT_0A(256'h07E0F83F07C0F83E07C1F03E0FC1F07E0F83F07C0F83E07C1F03E0F81F07C0F8),
    .INIT_0B(256'h81F07E0F81F07E0F81F07C0F83F07C0F83F07C1F83E07C1F83E0FC1F03E0F81F),
    .INIT_0C(256'h83F07C0F83F07E0F81F07E0F81F07E0F81F07E0F81F07E0F81F07E0F81F07E0F),
    .INIT_0D(256'h0F81F07E0FC1F03E07C1F83F07C0F81F07E0F81F03E0FC1F03E07C1F83E07C0F),
    .INIT_0E(256'hF03E07C0F81F07E0FC1F83F07C0F81F03E0FC1F83F07C0F81F03E0FC1F83E07C),
    .INIT_0F(256'h1F03E07C0F81F03E07C0F81F03E07C0F83F07E0FC1F83F07E0FC1F83F07C0F81),
    .INIT_10(256'h0F81F03E07E0FC1F83F07E07C0F81F03E07C0FC1F83F07E0FC1F83F07E0FC1F8),
    .INIT_11(256'h3E07E0FC0F81F83F07E07C0F81F83F07E07C0F81F83F07E07C0F81F83F07E0FC),
    .INIT_12(256'hE07C0FC1F81F03F07E07C0FC0F81F83F03E07E0FC0F81F03F07E07C0FC1F81F0),
    .INIT_13(256'h7C0FC0F81F81F03F03F07E07E0FC0F81F81F03F03E07E07C0FC1F81F83F03E07),
    .INIT_14(256'h7E0FC0FC0FC0F81F81F81F03F03F07E07E07E0FC0FC0F81F81F83F03F07E07E0),
    .INIT_15(256'hE07E07E07E07E07C0FC0FC0FC0FC0FC1F81F81F81F81F03F03F03F03E07E07E0),
    .INIT_16(256'h3F03F03F03F03F03F03F03F03F03F03F03F03F03F03F03F03F03F03F07E07E07),
    .INIT_17(256'h1F81F81F81FC0FC0FC0FC0FC0FE07E07E07E07E07E07E07F03F03F03F03F03F0),
    .INIT_18(256'hFC0FC0FC07E07E07F03F03F01F81F81FC0FC0FC0FE07E07E07F03F03F03F03F8),
    .INIT_19(256'h0FC07E07F03F01F81F80FC0FE07E03F03F01F81FC0FC0FE07E07F03F03F81F81),
    .INIT_1A(256'h0FC07E03F01F80FC0FE07F03F01F80FC07E07F03F01F80FC0FE07E03F01F81FC),
    .INIT_1B(256'hFC0FE07F03F80FC07E03F01F80FE07F03F81FC0FE07F03F81FC0FE07F03F81F8),
    .INIT_1C(256'h3F81FC07F03F80FC07F03F80FC07F03F80FC07F03F80FC07F03F81FC07E03F01),
    .INIT_1D(256'hFC07F01FC07F03F80FE03F81FC07F01FC0FE03F81FC07F01F80FE03F01FC07E0),
    .INIT_1E(256'h07F01FC07F01FC07F01FC07F01FC07F01FC07F01FC07F01FC0FE03F80FE03F80),
    .INIT_1F(256'h07F00FE03F80FF01FC07F01FC03F80FE03F80FE03FC07F01FC07F01FC07F01FC),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_032768_000 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n2734,open_n2735,open_n2736,open_n2737,open_n2738,open_n2739,open_n2740,1'b0,open_n2741}),
    .rsta(rsta),
    .doa({open_n2756,open_n2757,open_n2758,open_n2759,open_n2760,open_n2761,open_n2762,open_n2763,inst_doa_i4_000}));
  // address_offset=32768;data_offset=1;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h7FE007FE003FF003FF003FF001FF801FF801FFC00FFC00FFC007FE007FE007FF),
    .INIT_01(256'hC00FFC00FFE007FE007FE003FF003FF003FF801FF801FF800FFC00FFC00FFE00),
    .INIT_02(256'h1FF801FF800FFC00FFC00FFE007FE007FE003FF003FF003FF801FF801FF800FF),
    .INIT_03(256'hE007FF003FF003FF001FF801FF800FFC00FFC00FFE007FE007FF003FF003FF00),
    .INIT_04(256'h1FF801FFC00FFC00FFE007FE007FF003FF003FF801FF801FFC00FFC00FFE007F),
    .INIT_05(256'hC00FFC007FE007FE003FF003FF801FF801FFC00FFC007FE007FE003FF003FF00),
    .INIT_06(256'hFFC00FFE007FE003FF003FF801FF800FFC00FFE007FE003FF003FF801FF801FF),
    .INIT_07(256'h01FF800FFC007FE007FF003FF001FF800FFC00FFE007FE003FF003FF801FF800),
    .INIT_08(256'hE007FF003FF001FF800FFC007FE007FF003FF801FF800FFC007FE007FF003FF8),
    .INIT_09(256'hFE003FF001FF800FFC007FE003FF001FF800FFC007FE003FF003FF801FFC00FF),
    .INIT_0A(256'hFFE007FF003FF801FFC00FFE003FF001FF800FFC007FE003FF001FF800FFC007),
    .INIT_0B(256'h7FF001FF800FFE007FF003FF800FFC007FF003FF801FFC007FE003FF001FF800),
    .INIT_0C(256'h7FF003FF800FFE007FF001FF800FFE007FF001FF800FFE007FF001FF800FFE00),
    .INIT_0D(256'hFF800FFE003FF001FFC007FF003FF800FFE007FF001FFC00FFE003FF801FFC00),
    .INIT_0E(256'hF001FFC007FF001FFC007FF003FF800FFE003FF800FFC007FF001FFC007FE003),
    .INIT_0F(256'h00FFE003FF800FFE003FF800FFE003FF800FFE003FF800FFE003FF800FFC007F),
    .INIT_10(256'hFF800FFE001FFC007FF001FFC007FF001FFC003FF800FFE003FF800FFE003FF8),
    .INIT_11(256'h01FFE003FF8007FF001FFC007FF800FFE003FF8007FF001FFC007FF800FFE003),
    .INIT_12(256'hE003FFC007FF000FFE003FFC007FF800FFE001FFC007FF000FFE003FFC007FF0),
    .INIT_13(256'hFC003FF8007FF000FFF001FFE003FF8007FF000FFE001FFC003FF8007FF001FF),
    .INIT_14(256'hFE003FFC003FF8007FF800FFF000FFE001FFE003FFC007FF8007FF000FFE001F),
    .INIT_15(256'hE001FFE001FFE003FFC003FFC003FFC007FF8007FF800FFF000FFF001FFE001F),
    .INIT_16(256'h00FFF000FFF000FFF000FFF000FFF000FFF000FFF000FFF000FFF000FFE001FF),
    .INIT_17(256'hFF8007FF8003FFC003FFC003FFE001FFE001FFE001FFE000FFF000FFF000FFF0),
    .INIT_18(256'h03FFC003FFE001FFF000FFF0007FF8003FFC003FFE001FFE000FFF000FFF0007),
    .INIT_19(256'h003FFE000FFF0007FF8003FFE001FFF000FFF8003FFC001FFE000FFF0007FF80),
    .INIT_1A(256'h003FFE000FFF8003FFE000FFF0007FFC001FFF000FFF8003FFE001FFF0007FFC),
    .INIT_1B(256'h03FFE000FFF8003FFE000FFF8001FFF0007FFC001FFF0007FFC001FFF0007FF8),
    .INIT_1C(256'hFF8003FFF0007FFC000FFF8003FFF0007FFC000FFF8003FFF0007FFC001FFF00),
    .INIT_1D(256'h03FFF0003FFF0007FFE0007FFC000FFFC001FFF8003FFF0007FFE000FFFC001F),
    .INIT_1E(256'h000FFFC000FFFC000FFFC000FFFC000FFFC000FFFC000FFFC001FFF8001FFF80),
    .INIT_1F(256'h000FFFE0007FFF0003FFF0003FFF8001FFF8001FFFC000FFFC000FFFC000FFFC),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_032768_001 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n2792,open_n2793,open_n2794,open_n2795,open_n2796,open_n2797,open_n2798,1'b0,open_n2799}),
    .rsta(rsta),
    .doa({open_n2814,open_n2815,open_n2816,open_n2817,open_n2818,open_n2819,open_n2820,open_n2821,inst_doa_i4_001}));
  // address_offset=32768;data_offset=2;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFE00001FFFFF00000FFFFF000007FFFF800003FFFFC00003FFFFE00001FFFFF),
    .INIT_01(256'h3FFFFC00001FFFFE00001FFFFF00000FFFFF800007FFFF800003FFFFC00001FF),
    .INIT_02(256'h0007FFFF800003FFFFC00001FFFFE00001FFFFF00000FFFFF800007FFFF80000),
    .INIT_03(256'hE00000FFFFF00000FFFFF800007FFFFC00003FFFFE00001FFFFF00000FFFFF00),
    .INIT_04(256'hFFF800003FFFFC00001FFFFE00000FFFFF000007FFFF800003FFFFC00001FFFF),
    .INIT_05(256'h3FFFFC00001FFFFE00000FFFFF800007FFFFC00003FFFFE00001FFFFF00000FF),
    .INIT_06(256'h003FFFFE00001FFFFF000007FFFF800003FFFFE00001FFFFF000007FFFF80000),
    .INIT_07(256'h00007FFFFC00001FFFFF00000FFFFF800003FFFFE00001FFFFF000007FFFF800),
    .INIT_08(256'hE00000FFFFF000007FFFFC00001FFFFF000007FFFF800003FFFFE00000FFFFF8),
    .INIT_09(256'hFE00000FFFFF800003FFFFE00000FFFFF800003FFFFE00000FFFFF800003FFFF),
    .INIT_0A(256'hFFE00000FFFFF800003FFFFE00000FFFFF800003FFFFE00000FFFFF800003FFF),
    .INIT_0B(256'hFFF000007FFFFE00000FFFFF800003FFFFF000007FFFFC00001FFFFF000007FF),
    .INIT_0C(256'hFFF000007FFFFE00000FFFFF800001FFFFF000007FFFFE00000FFFFF800001FF),
    .INIT_0D(256'hFF800001FFFFF000003FFFFF000007FFFFE00000FFFFFC00001FFFFF800003FF),
    .INIT_0E(256'hF000003FFFFF000003FFFFF000007FFFFE000007FFFFC00000FFFFFC00001FFF),
    .INIT_0F(256'h00001FFFFF800001FFFFF800001FFFFF800001FFFFF800001FFFFF800003FFFF),
    .INIT_10(256'h007FFFFE000003FFFFF000003FFFFF000003FFFFF800001FFFFF800001FFFFF8),
    .INIT_11(256'hFFFFE000007FFFFF000003FFFFF800001FFFFF800000FFFFFC000007FFFFE000),
    .INIT_12(256'hE000003FFFFF000001FFFFFC000007FFFFE000003FFFFF000001FFFFFC00000F),
    .INIT_13(256'h03FFFFF800000FFFFFF000001FFFFF800000FFFFFE000003FFFFF800000FFFFF),
    .INIT_14(256'hFE000003FFFFF8000007FFFFF000001FFFFFE000003FFFFF800000FFFFFE0000),
    .INIT_15(256'h1FFFFFE000001FFFFFC000003FFFFFC000007FFFFF800000FFFFFF000001FFFF),
    .INIT_16(256'h00000FFFFFF000000FFFFFF000000FFFFFF000000FFFFFF000000FFFFFE00000),
    .INIT_17(256'hFF8000007FFFFFC000003FFFFFE000001FFFFFE000001FFFFFF000000FFFFFF0),
    .INIT_18(256'hFFFFC000001FFFFFF000000FFFFFF8000003FFFFFE000001FFFFFF000000FFFF),
    .INIT_19(256'hFFFFFE000000FFFFFF8000001FFFFFF0000007FFFFFC000001FFFFFF0000007F),
    .INIT_1A(256'hFFFFFE0000007FFFFFE000000FFFFFFC000000FFFFFF8000001FFFFFF0000003),
    .INIT_1B(256'hFFFFE0000007FFFFFE0000007FFFFFF0000003FFFFFF0000003FFFFFF0000007),
    .INIT_1C(256'hFF8000000FFFFFFC0000007FFFFFF0000003FFFFFF8000000FFFFFFC000000FF),
    .INIT_1D(256'h00000FFFFFFF0000001FFFFFFC0000003FFFFFF8000000FFFFFFE0000003FFFF),
    .INIT_1E(256'hFFFFFFC0000003FFFFFFC0000003FFFFFFC0000003FFFFFFC0000007FFFFFF80),
    .INIT_1F(256'h0000001FFFFFFF0000000FFFFFFF80000007FFFFFFC0000003FFFFFFC0000003),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_032768_002 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n2850,open_n2851,open_n2852,open_n2853,open_n2854,open_n2855,open_n2856,1'b0,open_n2857}),
    .rsta(rsta),
    .doa({open_n2872,open_n2873,open_n2874,open_n2875,open_n2876,open_n2877,open_n2878,open_n2879,inst_doa_i4_002}));
  // address_offset=32768;data_offset=3;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFE0000000000FFFFFFFFFF00000000007FFFFFFFFFC0000000001FFFFFFFFFF),
    .INIT_01(256'hFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFF80000000003FFFFFFF),
    .INIT_02(256'hFFFFFFFF80000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000007FFFF),
    .INIT_03(256'h1FFFFFFFFFF00000000007FFFFFFFFFC0000000001FFFFFFFFFF0000000000FF),
    .INIT_04(256'h0007FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFFC000000000),
    .INIT_05(256'h000003FFFFFFFFFE00000000007FFFFFFFFFC0000000001FFFFFFFFFF0000000),
    .INIT_06(256'h00000001FFFFFFFFFF00000000007FFFFFFFFFE0000000000FFFFFFFFFF80000),
    .INIT_07(256'h0000000003FFFFFFFFFF00000000007FFFFFFFFFE0000000000FFFFFFFFFF800),
    .INIT_08(256'hE0000000000FFFFFFFFFFC0000000000FFFFFFFFFF80000000001FFFFFFFFFF8),
    .INIT_09(256'hFE00000000007FFFFFFFFFE00000000007FFFFFFFFFE00000000007FFFFFFFFF),
    .INIT_0A(256'hFFE00000000007FFFFFFFFFE00000000007FFFFFFFFFE00000000007FFFFFFFF),
    .INIT_0B(256'hFFF00000000001FFFFFFFFFF80000000000FFFFFFFFFFC0000000000FFFFFFFF),
    .INIT_0C(256'hFFF00000000001FFFFFFFFFF80000000000FFFFFFFFFFE00000000007FFFFFFF),
    .INIT_0D(256'hFF80000000000FFFFFFFFFFF00000000001FFFFFFFFFFC00000000007FFFFFFF),
    .INIT_0E(256'hF00000000000FFFFFFFFFFF00000000001FFFFFFFFFFC00000000003FFFFFFFF),
    .INIT_0F(256'h00000000007FFFFFFFFFF800000000007FFFFFFFFFF800000000007FFFFFFFFF),
    .INIT_10(256'h00000001FFFFFFFFFFF00000000000FFFFFFFFFFF800000000007FFFFFFFFFF8),
    .INIT_11(256'h00001FFFFFFFFFFF000000000007FFFFFFFFFF800000000003FFFFFFFFFFE000),
    .INIT_12(256'h1FFFFFFFFFFF000000000003FFFFFFFFFFE00000000000FFFFFFFFFFFC000000),
    .INIT_13(256'hFFFFFFF800000000000FFFFFFFFFFF800000000001FFFFFFFFFFF80000000000),
    .INIT_14(256'hFE000000000007FFFFFFFFFFF000000000001FFFFFFFFFFF800000000001FFFF),
    .INIT_15(256'h0000001FFFFFFFFFFFC000000000003FFFFFFFFFFF800000000000FFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFFF000000000000FFFFFFFFFFFF000000000000FFFFFFFFFFFE00000),
    .INIT_17(256'hFF8000000000003FFFFFFFFFFFE000000000001FFFFFFFFFFFF000000000000F),
    .INIT_18(256'h00003FFFFFFFFFFFF0000000000007FFFFFFFFFFFE000000000000FFFFFFFFFF),
    .INIT_19(256'hFFFFFE0000000000007FFFFFFFFFFFF0000000000003FFFFFFFFFFFF00000000),
    .INIT_1A(256'h000001FFFFFFFFFFFFE0000000000003FFFFFFFFFFFF8000000000000FFFFFFF),
    .INIT_1B(256'hFFFFE0000000000001FFFFFFFFFFFFF0000000000000FFFFFFFFFFFFF0000000),
    .INIT_1C(256'h007FFFFFFFFFFFFC0000000000000FFFFFFFFFFFFF80000000000003FFFFFFFF),
    .INIT_1D(256'h000000000000FFFFFFFFFFFFFC00000000000007FFFFFFFFFFFFE00000000000),
    .INIT_1E(256'hFFFFFFC00000000000003FFFFFFFFFFFFFC00000000000003FFFFFFFFFFFFF80),
    .INIT_1F(256'hFFFFFFFFFFFFFF000000000000007FFFFFFFFFFFFFC00000000000003FFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_032768_003 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n2908,open_n2909,open_n2910,open_n2911,open_n2912,open_n2913,open_n2914,1'b0,open_n2915}),
    .rsta(rsta),
    .doa({open_n2930,open_n2931,open_n2932,open_n2933,open_n2934,open_n2935,open_n2936,open_n2937,inst_doa_i4_003}));
  // address_offset=32768;data_offset=4;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h001FFFFFFFFFFFFFFFFFFFF000000000000000000003FFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFF800000000000000000),
    .INIT_02(256'h000000007FFFFFFFFFFFFFFFFFFFE000000000000000000007FFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFF000000000000000000003FFFFFFFFFFFFFFFFFFFF000000000000),
    .INIT_04(256'h00000000000003FFFFFFFFFFFFFFFFFFFF000000000000000000003FFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFE000000000000000000003FFFFFFFFFFFFFFFFFFFF0000000),
    .INIT_06(256'h000000000000000000FFFFFFFFFFFFFFFFFFFFE000000000000000000007FFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFF000000000000000000001FFFFFFFFFFFFFFFFFFFF800),
    .INIT_08(256'hE000000000000000000003FFFFFFFFFFFFFFFFFFFF8000000000000000000007),
    .INIT_09(256'h01FFFFFFFFFFFFFFFFFFFFE000000000000000000001FFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFE000000000000000000001FFFFFFFFFFFFFFFFFFFFE0000000000000000000),
    .INIT_0B(256'h000FFFFFFFFFFFFFFFFFFFFF8000000000000000000003FFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFF0000000000000000000007FFFFFFFFFFFFFFFFFFFFE000000000000000000),
    .INIT_0D(256'h007FFFFFFFFFFFFFFFFFFFFF0000000000000000000003FFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hF0000000000000000000000FFFFFFFFFFFFFFFFFFFFFC0000000000000000000),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFF80000000000000000000007FFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'h0000000000000000000FFFFFFFFFFFFFFFFFFFFFF80000000000000000000007),
    .INIT_11(256'hFFFFFFFFFFFFFFFF00000000000000000000007FFFFFFFFFFFFFFFFFFFFFE000),
    .INIT_12(256'h000000000000FFFFFFFFFFFFFFFFFFFFFFE00000000000000000000003FFFFFF),
    .INIT_13(256'hFFFFFFF800000000000000000000007FFFFFFFFFFFFFFFFFFFFFF80000000000),
    .INIT_14(256'h01FFFFFFFFFFFFFFFFFFFFFFF000000000000000000000007FFFFFFFFFFFFFFF),
    .INIT_15(256'h0000000000000000003FFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000),
    .INIT_16(256'hFFFFFFFFFFF000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFE00000),
    .INIT_17(256'h007FFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000FFFFFFFFFFFFF),
    .INIT_18(256'h00000000000000000FFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000),
    .INIT_19(256'hFFFFFE0000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFF00000000),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFE00000000000000000000000007FFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'h00001FFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000FFFFFFF),
    .INIT_1C(256'h0000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000),
    .INIT_1D(256'h00000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000),
    .INIT_1E(256'hFFFFFFC0000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFF80),
    .INIT_1F(256'hFFFFFFFFFFFFFF00000000000000000000000000003FFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_032768_004 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n2966,open_n2967,open_n2968,open_n2969,open_n2970,open_n2971,open_n2972,1'b0,open_n2973}),
    .rsta(rsta),
    .doa({open_n2988,open_n2989,open_n2990,open_n2991,open_n2992,open_n2993,open_n2994,open_n2995,inst_doa_i4_004}));
  // address_offset=32768;data_offset=5;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'h000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000),
    .INIT_03(256'hFFFFFFFFFFF00000000000000000000000000000000000000000FFFFFFFFFFFF),
    .INIT_04(256'h0000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'h0000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000007FF),
    .INIT_08(256'hE000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'h00000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'h001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000),
    .INIT_0C(256'hFFF0000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'h000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'h0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000),
    .INIT_10(256'h000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000),
    .INIT_13(256'hFFFFFFF80000000000000000000000000000000000000000000007FFFFFFFFFF),
    .INIT_14(256'h0000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000),
    .INIT_16(256'hFFFFFFFFFFF000000000000000000000000000000000000000000000001FFFFF),
    .INIT_17(256'h000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000),
    .INIT_19(256'hFFFFFE00000000000000000000000000000000000000000000000000FFFFFFFF),
    .INIT_1A(256'h0000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000),
    .INIT_1E(256'hFFFFFFC00000000000000000000000000000000000000000000000000000007F),
    .INIT_1F(256'h00000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_032768_005 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n3024,open_n3025,open_n3026,open_n3027,open_n3028,open_n3029,open_n3030,1'b0,open_n3031}),
    .rsta(rsta),
    .doa({open_n3046,open_n3047,open_n3048,open_n3049,open_n3050,open_n3051,open_n3052,open_n3053,inst_doa_i4_005}));
  // address_offset=32768;data_offset=6;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'h00000000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000000),
    .INIT_03(256'h00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000),
    .INIT_06(256'h000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000),
    .INIT_08(256'h1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000),
    .INIT_0B(256'h0000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFF0000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'h000000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000001FFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000),
    .INIT_13(256'h00000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000),
    .INIT_16(256'h00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000),
    .INIT_19(256'h000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'h00000000000000000000000000000000000000000000000000001FFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFC000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_032768_006 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n3082,open_n3083,open_n3084,open_n3085,open_n3086,open_n3087,open_n3088,1'b0,open_n3089}),
    .rsta(rsta),
    .doa({open_n3104,open_n3105,open_n3106,open_n3107,open_n3108,open_n3109,open_n3110,open_n3111,inst_doa_i4_006}));
  // address_offset=32768;data_offset=7;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'h00000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'h00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'h000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'h00000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'h000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'h0000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_032768_007 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n3140,open_n3141,open_n3142,open_n3143,open_n3144,open_n3145,open_n3146,1'b0,open_n3147}),
    .rsta(rsta),
    .doa({open_n3162,open_n3163,open_n3164,open_n3165,open_n3166,open_n3167,open_n3168,open_n3169,inst_doa_i4_007}));
  // address_offset=32768;data_offset=8;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'h000000000000000000000000000000000000000000000000000000000FFFFFFF),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'h0000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'h0000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_032768_008 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n3198,open_n3199,open_n3200,open_n3201,open_n3202,open_n3203,open_n3204,1'b0,open_n3205}),
    .rsta(rsta),
    .doa({open_n3220,open_n3221,open_n3222,open_n3223,open_n3224,open_n3225,open_n3226,open_n3227,inst_doa_i4_008}));
  // address_offset=32768;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'h000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_032768_009 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n3256,open_n3257,open_n3258,open_n3259,open_n3260,open_n3261,open_n3262,1'b0,open_n3263}),
    .rsta(rsta),
    .doa({open_n3278,open_n3279,open_n3280,open_n3281,open_n3282,open_n3283,open_n3284,open_n3285,inst_doa_i4_009}));
  // address_offset=32768;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'h0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_032768_010 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n3314,open_n3315,open_n3316,open_n3317,open_n3318,open_n3319,open_n3320,1'b0,open_n3321}),
    .rsta(rsta),
    .doa({open_n3336,open_n3337,open_n3338,open_n3339,open_n3340,open_n3341,open_n3342,open_n3343,inst_doa_i4_010}));
  // address_offset=32768;data_offset=11;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_032768_011 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n3372,open_n3373,open_n3374,open_n3375,open_n3376,open_n3377,open_n3378,1'b0,open_n3379}),
    .rsta(rsta),
    .doa({open_n3394,open_n3395,open_n3396,open_n3397,open_n3398,open_n3399,open_n3400,open_n3401,inst_doa_i4_011}));
  // address_offset=40960;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFC07F80FF01FC03F80FF01FC03F80FF01FC07F80FE01FC07F00FE03F80FF01FC),
    .INIT_01(256'hFF01FE01FC03F807F00FE01FC03F807F00FE01FC03F807F01FE03FC07F80FE01),
    .INIT_02(256'hE03FC03FC07F807F80FF00FF01FE01FC03FC07F807F00FF01FE01FC03F807F80),
    .INIT_03(256'hF807F807F807F807F807F807F807F807F807F807F00FF00FF00FF01FE01FE01F),
    .INIT_04(256'h807F807FC03FC03FE01FE01FE00FF00FF00FF00FF807F807F807F807F807F807),
    .INIT_05(256'hF007F803FC01FE00FF007F803FC01FE00FF00FF807F803FC03FE01FE00FF00FF),
    .INIT_06(256'h00FF803FE00FF007FC01FE00FF803FC01FF00FF803FC01FF00FF803FC01FE00F),
    .INIT_07(256'hE007FC01FF007FC01FF007FE00FF803FE00FF803FE01FF007FC01FF007FC01FF),
    .INIT_08(256'h01FF803FF007FE00FFC01FF803FE007FC01FF803FE007FC01FF003FE00FF803F),
    .INIT_09(256'h801FF801FF801FF803FF003FF003FE007FE00FFC00FF801FF803FF007FE00FFC),
    .INIT_0A(256'h07FE007FF003FF003FF801FF801FF801FF800FFC00FFC00FFC00FFC00FFC00FF),
    .INIT_0B(256'h01FFC007FF003FF800FFC007FF003FF801FFC007FE003FF003FF801FFC00FFC0),
    .INIT_0C(256'hFF8007FF001FFC003FF800FFE003FF800FFE003FF800FFE003FF800FFE003FF8),
    .INIT_0D(256'hFFC003FFC003FFC003FF8007FF800FFF000FFE001FFC003FF8007FF001FFE003),
    .INIT_0E(256'h003FFE001FFF000FFF0007FF8007FFC003FFC003FFC003FFE001FFE001FFE001),
    .INIT_0F(256'h00FFF8001FFF0007FFC001FFF0007FFC001FFF0007FF8003FFE000FFF0007FFC),
    .INIT_10(256'hF0003FFF0003FFF0003FFF0003FFE0007FFE000FFFC000FFF8001FFF0007FFE0),
    .INIT_11(256'h000FFFE0003FFF8000FFFC0007FFF0003FFF8000FFFC000FFFE0007FFE0003FF),
    .INIT_12(256'hC0003FFFC0003FFFC0003FFFC0003FFFC0007FFF8000FFFF0001FFFC0007FFF8),
    .INIT_13(256'h07FFFE0000FFFFC0001FFFF00007FFFC0001FFFE0000FFFF80007FFF80003FFF),
    .INIT_14(256'h03FFFF80000FFFFC00007FFFF00003FFFF00003FFFF80001FFFF00003FFFF000),
    .INIT_15(256'hC00001FFFFF000007FFFF800007FFFF800007FFFF800007FFFF00001FFFFE000),
    .INIT_16(256'h00007FFFFF000001FFFFF800001FFFFFC00000FFFFF800001FFFFF000007FFFF),
    .INIT_17(256'hF0000003FFFFFE000000FFFFFF8000003FFFFFE000001FFFFFE000003FFFFFC0),
    .INIT_18(256'h003FFFFFFE0000000FFFFFFF80000007FFFFFF8000000FFFFFFE0000007FFFFF),
    .INIT_19(256'h001FFFFFFFF800000001FFFFFFFE00000001FFFFFFFE00000003FFFFFFF00000),
    .INIT_1A(256'hF00000000007FFFFFFFFF0000000001FFFFFFFFF0000000007FFFFFFFF000000),
    .INIT_1B(256'h00000000FFFFFFFFFFFFC000000000007FFFFFFFFFFC00000000003FFFFFFFFF),
    .INIT_1C(256'h0000000000000001FFFFFFFFFFFFFFF800000000000003FFFFFFFFFFFFF80000),
    .INIT_1D(256'h1FFFFFFFFFFFFFFFFFFFFFFF800000000000000000001FFFFFFFFFFFFFFFFFF0),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000003FFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_040960_000 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n3430,open_n3431,open_n3432,open_n3433,open_n3434,open_n3435,open_n3436,1'b0,open_n3437}),
    .rsta(rsta),
    .doa({open_n3452,open_n3453,open_n3454,open_n3455,open_n3456,open_n3457,open_n3458,open_n3459,inst_doa_i5_000}));
  // address_offset=40960;data_offset=1;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h03FFF8000FFFC0007FFF0003FFF8000FFFC0007FFE0003FFF0001FFF8000FFFC),
    .INIT_01(256'hFF0001FFFC0007FFF0001FFFC0007FFF0001FFFC0007FFF0001FFFC0007FFE00),
    .INIT_02(256'h1FFFC0003FFF80007FFF0000FFFE0003FFFC0007FFF0000FFFE0003FFF80007F),
    .INIT_03(256'h07FFF80007FFF80007FFF80007FFF80007FFF8000FFFF0000FFFF0001FFFE000),
    .INIT_04(256'h7FFF80003FFFC0001FFFE0001FFFF0000FFFF00007FFF80007FFF80007FFF800),
    .INIT_05(256'hF00007FFFC0001FFFF00007FFFC0001FFFF00007FFF80003FFFE0001FFFF0000),
    .INIT_06(256'hFFFF80001FFFF00003FFFE00007FFFC0000FFFF80003FFFF00007FFFC0001FFF),
    .INIT_07(256'h1FFFFC0000FFFFC0000FFFFE00007FFFE00007FFFE0000FFFFC0000FFFFC0000),
    .INIT_08(256'hFFFF80000FFFFE00003FFFF80001FFFFC00007FFFE00003FFFF00001FFFF8000),
    .INIT_09(256'h800007FFFF800007FFFF00000FFFFE00001FFFFC00007FFFF80000FFFFE00003),
    .INIT_0A(256'hFFFE00000FFFFF000007FFFF800007FFFF800003FFFFC00003FFFFC00003FFFF),
    .INIT_0B(256'hFFFFC00000FFFFF800003FFFFF000007FFFFC00001FFFFF000007FFFFC00003F),
    .INIT_0C(256'hFF800000FFFFFC000007FFFFE000007FFFFE000007FFFFE000007FFFFE000007),
    .INIT_0D(256'h003FFFFFC000003FFFFF8000007FFFFF000001FFFFFC000007FFFFF000001FFF),
    .INIT_0E(256'h000001FFFFFF000000FFFFFF8000003FFFFFC000003FFFFFE000001FFFFFE000),
    .INIT_0F(256'h000007FFFFFF0000003FFFFFF0000003FFFFFF0000007FFFFFE000000FFFFFFC),
    .INIT_10(256'h0FFFFFFF0000000FFFFFFF0000001FFFFFFE0000003FFFFFF8000000FFFFFFE0),
    .INIT_11(256'h0000001FFFFFFF80000003FFFFFFF00000007FFFFFFC0000001FFFFFFE000000),
    .INIT_12(256'hC00000003FFFFFFFC00000003FFFFFFFC00000007FFFFFFF00000003FFFFFFF8),
    .INIT_13(256'h000001FFFFFFFFC00000000FFFFFFFFC00000001FFFFFFFF800000007FFFFFFF),
    .INIT_14(256'hFFFFFF8000000003FFFFFFFFF000000000FFFFFFFFF800000000FFFFFFFFF000),
    .INIT_15(256'h3FFFFFFFFFF00000000007FFFFFFFFF80000000007FFFFFFFFF0000000001FFF),
    .INIT_16(256'hFFFFFFFFFF000000000007FFFFFFFFFFC00000000007FFFFFFFFFF0000000000),
    .INIT_17(256'hF0000000000001FFFFFFFFFFFF8000000000001FFFFFFFFFFFE000000000003F),
    .INIT_18(256'hFFFFFFFFFE000000000000007FFFFFFFFFFFFF80000000000001FFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFF80000000000000001FFFFFFFFFFFFFFFE000000000000000FFFFF),
    .INIT_1A(256'hF00000000000000000000FFFFFFFFFFFFFFFFFFF000000000000000000FFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFC00000000000000000000003FFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000007FFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000F),
    .INIT_1E(256'h000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_040960_001 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n3488,open_n3489,open_n3490,open_n3491,open_n3492,open_n3493,open_n3494,1'b0,open_n3495}),
    .rsta(rsta),
    .doa({open_n3510,open_n3511,open_n3512,open_n3513,open_n3514,open_n3515,open_n3516,open_n3517,inst_doa_i5_001}));
  // address_offset=40960;data_offset=2;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFF80000003FFFFFFF00000007FFFFFFC0000001FFFFFFF00000007FFFFFFC),
    .INIT_01(256'h00FFFFFFFC0000000FFFFFFFC0000000FFFFFFFC0000000FFFFFFFC0000001FF),
    .INIT_02(256'h00003FFFFFFF80000000FFFFFFFE00000003FFFFFFF00000001FFFFFFF800000),
    .INIT_03(256'h000007FFFFFFF800000007FFFFFFF800000007FFFFFFF00000000FFFFFFFE000),
    .INIT_04(256'h00007FFFFFFFC00000001FFFFFFFF00000000FFFFFFFF800000007FFFFFFF800),
    .INIT_05(256'h0FFFFFFFFC00000000FFFFFFFFC00000000FFFFFFFF800000001FFFFFFFF0000),
    .INIT_06(256'hFFFF800000000FFFFFFFFE000000003FFFFFFFF800000000FFFFFFFFC0000000),
    .INIT_07(256'h000003FFFFFFFFC000000001FFFFFFFFE000000001FFFFFFFFC000000003FFFF),
    .INIT_08(256'hFFFF8000000001FFFFFFFFF8000000003FFFFFFFFE000000000FFFFFFFFF8000),
    .INIT_09(256'h7FFFFFFFFF8000000000FFFFFFFFFE0000000003FFFFFFFFF8000000001FFFFF),
    .INIT_0A(256'h0001FFFFFFFFFF00000000007FFFFFFFFF80000000003FFFFFFFFFC000000000),
    .INIT_0B(256'h00003FFFFFFFFFF80000000000FFFFFFFFFFC0000000000FFFFFFFFFFC000000),
    .INIT_0C(256'h007FFFFFFFFFFC00000000001FFFFFFFFFFE00000000001FFFFFFFFFFE000000),
    .INIT_0D(256'hFFFFFFFFC000000000007FFFFFFFFFFF000000000003FFFFFFFFFFF000000000),
    .INIT_0E(256'h000000000000FFFFFFFFFFFF8000000000003FFFFFFFFFFFE000000000001FFF),
    .INIT_0F(256'hFFFFFFFFFFFF0000000000000FFFFFFFFFFFFF0000000000001FFFFFFFFFFFFC),
    .INIT_10(256'h00000000FFFFFFFFFFFFFF00000000000001FFFFFFFFFFFFF80000000000001F),
    .INIT_11(256'h000000000000007FFFFFFFFFFFFFF000000000000003FFFFFFFFFFFFFE000000),
    .INIT_12(256'hC0000000000000003FFFFFFFFFFFFFFFC000000000000000FFFFFFFFFFFFFFF8),
    .INIT_13(256'h000000000000003FFFFFFFFFFFFFFFFC00000000000000007FFFFFFFFFFFFFFF),
    .INIT_14(256'h0000007FFFFFFFFFFFFFFFFFF0000000000000000007FFFFFFFFFFFFFFFFF000),
    .INIT_15(256'hFFFFFFFFFFF000000000000000000007FFFFFFFFFFFFFFFFFFF0000000000000),
    .INIT_16(256'h0000000000FFFFFFFFFFFFFFFFFFFFFFC000000000000000000000FFFFFFFFFF),
    .INIT_17(256'hF00000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFE0000000000000),
    .INIT_18(256'hFFFFFFFFFE00000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFF800000000000000000000000000000001FFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hF000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'h000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_040960_002 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n3546,open_n3547,open_n3548,open_n3549,open_n3550,open_n3551,open_n3552,1'b0,open_n3553}),
    .rsta(rsta),
    .doa({open_n3568,open_n3569,open_n3570,open_n3571,open_n3572,open_n3573,open_n3574,open_n3575,inst_doa_i5_002}));
  // address_offset=40960;data_offset=3;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h000007FFFFFFFFFFFFFF000000000000003FFFFFFFFFFFFFF000000000000003),
    .INIT_01(256'h0000000003FFFFFFFFFFFFFFC000000000000003FFFFFFFFFFFFFFC000000000),
    .INIT_02(256'h0000000000007FFFFFFFFFFFFFFE000000000000000FFFFFFFFFFFFFFF800000),
    .INIT_03(256'h00000000000007FFFFFFFFFFFFFFF8000000000000000FFFFFFFFFFFFFFFE000),
    .INIT_04(256'h0000000000003FFFFFFFFFFFFFFFF00000000000000007FFFFFFFFFFFFFFF800),
    .INIT_05(256'h0000000003FFFFFFFFFFFFFFFFC00000000000000007FFFFFFFFFFFFFFFF0000),
    .INIT_06(256'h00007FFFFFFFFFFFFFFFFE000000000000000007FFFFFFFFFFFFFFFFC0000000),
    .INIT_07(256'hFFFFFFFFFFFFFFC000000000000000001FFFFFFFFFFFFFFFFFC0000000000000),
    .INIT_08(256'hFFFF80000000000000000007FFFFFFFFFFFFFFFFFE0000000000000000007FFF),
    .INIT_09(256'h00000000007FFFFFFFFFFFFFFFFFFE00000000000000000007FFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFF000000000000000000007FFFFFFFFFFFFFFFFFFFC000000000),
    .INIT_0B(256'h0000000000000007FFFFFFFFFFFFFFFFFFFFC000000000000000000003FFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFC0000000000000000000001FFFFFFFFFFFFFFFFFFFFFE000000),
    .INIT_0D(256'h000000003FFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000FFFFFFFFF),
    .INIT_0E(256'h0000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFE000000000000000),
    .INIT_0F(256'hFFFFFFFFFFFF00000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFC),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000007FFFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000001FFFFFF),
    .INIT_12(256'h3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000007),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000FFF),
    .INIT_15(256'hFFFFFFFFFFF0000000000000000000000000000000000000000FFFFFFFFFFFFF),
    .INIT_16(256'h000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'h0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000),
    .INIT_18(256'hFFFFFFFFFE000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hF000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'h00000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_040960_003 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n3604,open_n3605,open_n3606,open_n3607,open_n3608,open_n3609,open_n3610,1'b0,open_n3611}),
    .rsta(rsta),
    .doa({open_n3626,open_n3627,open_n3628,open_n3629,open_n3630,open_n3631,open_n3632,open_n3633,inst_doa_i5_003}));
  // address_offset=40960;data_offset=4;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000FFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000003FFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000007FFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000001FFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000007FF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000FFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000003FFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFC000000000000000000000000000000000003FFFFFFFFFFFFF),
    .INIT_08(256'hFFFF80000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'h000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'h00000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000),
    .INIT_0C(256'hFFFFFFFFFFFFFC00000000000000000000000000000000000000000001FFFFFF),
    .INIT_0D(256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000),
    .INIT_0F(256'hFFFFFFFFFFFF0000000000000000000000000000000000000000000000000003),
    .INIT_10(256'h0000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000),
    .INIT_12(256'h000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFFF00000000000000000000000000000000000000000000000000000),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'h000000000000000000000000000000000000000000000000001FFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFE000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'h0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_040960_004 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n3662,open_n3663,open_n3664,open_n3665,open_n3666,open_n3667,open_n3668,1'b0,open_n3669}),
    .rsta(rsta),
    .doa({open_n3684,open_n3685,open_n3686,open_n3687,open_n3688,open_n3689,open_n3690,open_n3691,inst_doa_i5_004}));
  // address_offset=40960;data_offset=5;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000),
    .INIT_03(256'h000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000),
    .INIT_05(256'h000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000),
    .INIT_07(256'h000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFF800000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000003FFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000),
    .INIT_0C(256'h00000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000),
    .INIT_0F(256'h000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'h00000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'hFFFFFFFFFFF00000000000000000000000000000000000000000000000000000),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'h0000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_040960_005 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n3720,open_n3721,open_n3722,open_n3723,open_n3724,open_n3725,open_n3726,1'b0,open_n3727}),
    .rsta(rsta),
    .doa({open_n3742,open_n3743,open_n3744,open_n3745,open_n3746,open_n3747,open_n3748,open_n3749,inst_doa_i5_005}));
  // address_offset=40960;data_offset=6;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'h00000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000000000),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'h00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000001FFFFFFFFFFFFFFF),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'h00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_040960_006 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n3778,open_n3779,open_n3780,open_n3781,open_n3782,open_n3783,open_n3784,1'b0,open_n3785}),
    .rsta(rsta),
    .doa({open_n3800,open_n3801,open_n3802,open_n3803,open_n3804,open_n3805,open_n3806,open_n3807,inst_doa_i5_006}));
  // address_offset=40960;data_offset=7;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'h0000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h00000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_040960_007 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n3836,open_n3837,open_n3838,open_n3839,open_n3840,open_n3841,open_n3842,1'b0,open_n3843}),
    .rsta(rsta),
    .doa({open_n3858,open_n3859,open_n3860,open_n3861,open_n3862,open_n3863,open_n3864,open_n3865,inst_doa_i5_007}));
  // address_offset=40960;data_offset=8;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'h0000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_040960_008 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n3894,open_n3895,open_n3896,open_n3897,open_n3898,open_n3899,open_n3900,1'b0,open_n3901}),
    .rsta(rsta),
    .doa({open_n3916,open_n3917,open_n3918,open_n3919,open_n3920,open_n3921,open_n3922,open_n3923,inst_doa_i5_008}));
  // address_offset=40960;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'h0000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_040960_009 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n3952,open_n3953,open_n3954,open_n3955,open_n3956,open_n3957,open_n3958,1'b0,open_n3959}),
    .rsta(rsta),
    .doa({open_n3974,open_n3975,open_n3976,open_n3977,open_n3978,open_n3979,open_n3980,open_n3981,inst_doa_i5_009}));
  // address_offset=40960;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_040960_010 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n4010,open_n4011,open_n4012,open_n4013,open_n4014,open_n4015,open_n4016,1'b0,open_n4017}),
    .rsta(rsta),
    .doa({open_n4032,open_n4033,open_n4034,open_n4035,open_n4036,open_n4037,open_n4038,open_n4039,inst_doa_i5_010}));
  // address_offset=49152;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFF8000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'h1FFFFFFFFFFFFFFFFFF000000000000000000003FFFFFFFFFFFFFFFFFFFFFFF0),
    .INIT_03(256'h00003FFFFFFFFFFFFF800000000000003FFFFFFFFFFFFFFF0000000000000000),
    .INIT_04(256'hFFFFFFFFF800000000007FFFFFFFFFFC000000000007FFFFFFFFFFFE00000000),
    .INIT_05(256'h000001FFFFFFFFC000000001FFFFFFFFF0000000001FFFFFFFFFC0000000001F),
    .INIT_06(256'h00001FFFFFFF80000000FFFFFFFF00000000FFFFFFFF000000003FFFFFFFF000),
    .INIT_07(256'hFFFFFC000000FFFFFFE0000003FFFFFFC0000003FFFFFFE0000000FFFFFFF800),
    .INIT_08(256'h07FFFFF800000FFFFFF000000FFFFFF8000003FFFFFE000000FFFFFF8000001F),
    .INIT_09(256'hFFFFC00001FFFFF000003FFFFE000007FFFFF000003FFFFF000001FFFFFC0000),
    .INIT_0A(256'h000FFFFF00001FFFFC00003FFFFC00003FFFFC00003FFFFC00001FFFFF000007),
    .INIT_0B(256'h001FFFF80001FFFF00003FFFF80001FFFF80001FFFFC00007FFFE00003FFFF80),
    .INIT_0C(256'hFFF80003FFFC0003FFFE0000FFFF00007FFFC0001FFFF00003FFFE0000FFFFC0),
    .INIT_0D(256'h3FFFC0007FFF0001FFFE0003FFFC0007FFF80007FFF80007FFF80007FFF80007),
    .INIT_0E(256'hFF8000FFFC000FFFE0007FFE0003FFF8001FFFC0007FFE0003FFF8000FFFE000),
    .INIT_0F(256'h0FFFC001FFF0003FFE0007FFE000FFFC000FFF8001FFF8001FFF8001FFF8001F),
    .INIT_10(256'h7FFC001FFE000FFF8003FFC001FFF0007FFC001FFF0007FFC001FFF0003FFE00),
    .INIT_11(256'h000FFF000FFF000FFF8007FF8007FF8007FFC003FFC001FFE001FFF000FFF800),
    .INIT_12(256'h800FFF001FFC003FF8007FF000FFE001FFE003FFC003FF8007FF8007FF8007FF),
    .INIT_13(256'h3FF800FFE003FF800FFE003FF800FFE003FF800FFE003FF8007FF001FFC003FF),
    .INIT_14(256'h07FE007FF003FF801FF800FFC007FF003FF801FFC007FE003FF801FFC007FF00),
    .INIT_15(256'hFE007FE007FE007FE007FE007FE003FF003FF003FF003FF801FF801FFC00FFC0),
    .INIT_16(256'h7FE00FFC01FF803FF003FE007FE00FFC00FF801FF801FF803FF003FF003FF003),
    .INIT_17(256'hF803FE00FF801FF007FC00FF803FF007FC00FF803FF007FE00FFC01FF803FF00),
    .INIT_18(256'hFF007FC01FF007FC01FF00FF803FE00FF803FE00FFC01FF007FC01FF007FC00F),
    .INIT_19(256'hE00FF007FC03FE01FF007F803FE01FF007F803FE00FF007FC01FE00FF803FE01),
    .INIT_1A(256'hFE01FE00FF00FF807F803FC03FE01FE00FF007F803FC01FE00FF007F803FC01F),
    .INIT_1B(256'hC03FC03FC03FC03FC03FC03FE01FE01FE01FE00FF00FF00FF807F807FC03FC03),
    .INIT_1C(256'hF00FF00FF01FE01FE01FE01FC03FC03FC03FC03FC03FC03FC03FC03FC03FC03F),
    .INIT_1D(256'h03FC03F807F00FF01FE01FC03FC07F807F00FF01FE01FE03FC03FC07F807F80F),
    .INIT_1E(256'h00FE03FC07F80FF01FC03F807F00FE01FC03F807F00FE01FC03F807F00FF01FE),
    .INIT_1F(256'h7F01FE03F80FE01FC07F00FE03FC07F01FE03F807F01FE03F807F01FE03FC07F),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_049152_000 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n4068,open_n4069,open_n4070,open_n4071,open_n4072,open_n4073,open_n4074,1'b0,open_n4075}),
    .rsta(rsta),
    .doa({open_n4090,open_n4091,open_n4092,open_n4093,open_n4094,open_n4095,open_n4096,open_n4097,inst_doa_i6_000}));
  // address_offset=49152;data_offset=1;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000),
    .INIT_02(256'hE000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFC0000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFF800000000000000000000007FFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFE000000000000000001FFFFFFFFFFFFFFFFFFE00000000000000000001F),
    .INIT_06(256'hFFFFE000000000000000FFFFFFFFFFFFFFFF00000000000000003FFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFF00000000000003FFFFFFFFFFFFFC00000000000000FFFFFFFFFF),
    .INIT_08(256'hF800000000000FFFFFFFFFFFF0000000000003FFFFFFFFFFFF0000000000001F),
    .INIT_09(256'h0000000001FFFFFFFFFFC00000000007FFFFFFFFFFC00000000001FFFFFFFFFF),
    .INIT_0A(256'hFFF0000000001FFFFFFFFFC0000000003FFFFFFFFFC0000000001FFFFFFFFFF8),
    .INIT_0B(256'h001FFFFFFFFE000000003FFFFFFFFE000000001FFFFFFFFF8000000003FFFFFF),
    .INIT_0C(256'hFFFFFFFC00000003FFFFFFFF000000007FFFFFFFE000000003FFFFFFFF000000),
    .INIT_0D(256'h3FFFFFFF80000001FFFFFFFC00000007FFFFFFF800000007FFFFFFF800000007),
    .INIT_0E(256'h000000FFFFFFF00000007FFFFFFC0000001FFFFFFF80000003FFFFFFF0000000),
    .INIT_0F(256'h0FFFFFFE0000003FFFFFF8000000FFFFFFF0000001FFFFFFE0000001FFFFFFE0),
    .INIT_10(256'h7FFFFFE000000FFFFFFC000001FFFFFF8000001FFFFFF8000001FFFFFFC00000),
    .INIT_11(256'h000FFFFFF000000FFFFFF8000007FFFFF8000003FFFFFE000001FFFFFF000000),
    .INIT_12(256'hFFF000001FFFFFC000007FFFFF000001FFFFFC000003FFFFF8000007FFFFF800),
    .INIT_13(256'hC00000FFFFFC00000FFFFFC00000FFFFFC00000FFFFFC000007FFFFE000003FF),
    .INIT_14(256'hF800007FFFFC00001FFFFF000007FFFFC00001FFFFF800003FFFFE000007FFFF),
    .INIT_15(256'hFFFF800007FFFF800007FFFF800003FFFFC00003FFFFC00001FFFFE00000FFFF),
    .INIT_16(256'h80000FFFFE00003FFFFC00007FFFF00000FFFFE00001FFFFC00003FFFFC00003),
    .INIT_17(256'h0003FFFF00001FFFF80000FFFFC00007FFFF00003FFFF80000FFFFE00003FFFF),
    .INIT_18(256'h00007FFFE00007FFFE0000FFFFC0000FFFFC0000FFFFE00007FFFE00007FFFF0),
    .INIT_19(256'hFFF00007FFFC0001FFFF80003FFFE00007FFFC0000FFFF80001FFFF00003FFFE),
    .INIT_1A(256'h0001FFFF0000FFFF80003FFFC0001FFFF00007FFFC0001FFFF00007FFFC0001F),
    .INIT_1B(256'h003FFFC0003FFFC0003FFFC0001FFFE0001FFFF0000FFFF00007FFF80003FFFC),
    .INIT_1C(256'h000FFFF0001FFFE0001FFFE0003FFFC0003FFFC0003FFFC0003FFFC0003FFFC0),
    .INIT_1D(256'hFC0003FFF8000FFFE0001FFFC0007FFF8000FFFE0001FFFC0003FFF80007FFF0),
    .INIT_1E(256'h00FFFC0007FFF0001FFFC0007FFF0001FFFC0007FFF0001FFFC0007FFF0001FF),
    .INIT_1F(256'h7FFE0003FFF0001FFF8000FFFC0007FFE0003FFF8001FFFC0007FFE0003FFF80),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_049152_001 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n4126,open_n4127,open_n4128,open_n4129,open_n4130,open_n4131,open_n4132,1'b0,open_n4133}),
    .rsta(rsta),
    .doa({open_n4148,open_n4149,open_n4150,open_n4151,open_n4152,open_n4153,open_n4154,open_n4155,inst_doa_i6_001}));
  // address_offset=49152;data_offset=2;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000),
    .INIT_03(256'h000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000001F),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000003FFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000FFFFFFFFFF),
    .INIT_08(256'h0000000000000FFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000001F),
    .INIT_09(256'hFFFFFFFFFE0000000000000000000007FFFFFFFFFFFFFFFFFFFFFE0000000000),
    .INIT_0A(256'h0000000000001FFFFFFFFFFFFFFFFFFFC00000000000000000001FFFFFFFFFFF),
    .INIT_0B(256'h001FFFFFFFFFFFFFFFFFC000000000000000001FFFFFFFFFFFFFFFFFFC000000),
    .INIT_0C(256'hFFFFFFFFFFFFFFFC00000000000000007FFFFFFFFFFFFFFFFC00000000000000),
    .INIT_0D(256'h3FFFFFFFFFFFFFFE0000000000000007FFFFFFFFFFFFFFF80000000000000007),
    .INIT_0E(256'h000000FFFFFFFFFFFFFF800000000000001FFFFFFFFFFFFFFC00000000000000),
    .INIT_0F(256'hF00000000000003FFFFFFFFFFFFF00000000000001FFFFFFFFFFFFFE00000000),
    .INIT_10(256'h7FFFFFFFFFFFF0000000000001FFFFFFFFFFFFE0000000000001FFFFFFFFFFFF),
    .INIT_11(256'hFFF000000000000FFFFFFFFFFFF8000000000003FFFFFFFFFFFE000000000000),
    .INIT_12(256'h000000001FFFFFFFFFFF800000000001FFFFFFFFFFFC000000000007FFFFFFFF),
    .INIT_13(256'h000000FFFFFFFFFFF00000000000FFFFFFFFFFF000000000007FFFFFFFFFFC00),
    .INIT_14(256'h0000007FFFFFFFFFE00000000007FFFFFFFFFE00000000003FFFFFFFFFF80000),
    .INIT_15(256'h0000000007FFFFFFFFF80000000003FFFFFFFFFC0000000001FFFFFFFFFF0000),
    .INIT_16(256'hFFFFF0000000003FFFFFFFFF8000000000FFFFFFFFFE0000000003FFFFFFFFFC),
    .INIT_17(256'h0003FFFFFFFFE000000000FFFFFFFFF8000000003FFFFFFFFF0000000003FFFF),
    .INIT_18(256'hFFFF8000000007FFFFFFFF000000000FFFFFFFFF0000000007FFFFFFFF800000),
    .INIT_19(256'h00000007FFFFFFFE000000003FFFFFFFF800000000FFFFFFFFE000000003FFFF),
    .INIT_1A(256'h0001FFFFFFFF000000003FFFFFFFE000000007FFFFFFFE000000007FFFFFFFE0),
    .INIT_1B(256'h003FFFFFFFC00000003FFFFFFFE00000001FFFFFFFF000000007FFFFFFFC0000),
    .INIT_1C(256'h000FFFFFFFE00000001FFFFFFFC00000003FFFFFFFC00000003FFFFFFFC00000),
    .INIT_1D(256'h000003FFFFFFF00000001FFFFFFF80000000FFFFFFFE00000003FFFFFFF80000),
    .INIT_1E(256'hFF00000007FFFFFFE00000007FFFFFFE00000007FFFFFFE00000007FFFFFFE00),
    .INIT_1F(256'h7FFFFFFC0000001FFFFFFF00000007FFFFFFC0000001FFFFFFF80000003FFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_049152_002 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n4184,open_n4185,open_n4186,open_n4187,open_n4188,open_n4189,open_n4190,1'b0,open_n4191}),
    .rsta(rsta),
    .doa({open_n4206,open_n4207,open_n4208,open_n4209,open_n4210,open_n4211,open_n4212,open_n4213,inst_doa_i6_002}));
  // address_offset=49152;data_offset=3;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000000000000000000000000),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'h000000000000000000000000000000000000000000000000000000000000001F),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000),
    .INIT_07(256'h000000000000000000000000000000000000000000000000000000FFFFFFFFFF),
    .INIT_08(256'h0000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000),
    .INIT_0A(256'hFFFFFFFFFFFFE0000000000000000000000000000000000000001FFFFFFFFFFF),
    .INIT_0B(256'hFFE000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'h000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hC0000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8),
    .INIT_0E(256'hFFFFFF00000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFFFFFFC000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'h7FFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000001FFFFFFFFFFFF),
    .INIT_11(256'h000000000000000FFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000),
    .INIT_12(256'hFFFFFFFFE00000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF800000000),
    .INIT_13(256'h000000FFFFFFFFFFFFFFFFFFFFFF00000000000000000000007FFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFF8000000000000000000007FFFFFFFFFFFFFFFFFFFFC000000000000000),
    .INIT_15(256'h0000000007FFFFFFFFFFFFFFFFFFFC00000000000000000001FFFFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFFFFFFC0000000000000000000FFFFFFFFFFFFFFFFFFFC0000000000),
    .INIT_17(256'hFFFC000000000000000000FFFFFFFFFFFFFFFFFFC0000000000000000003FFFF),
    .INIT_18(256'h00000000000007FFFFFFFFFFFFFFFFF0000000000000000007FFFFFFFFFFFFFF),
    .INIT_19(256'h00000007FFFFFFFFFFFFFFFFC00000000000000000FFFFFFFFFFFFFFFFFC0000),
    .INIT_1A(256'h0001FFFFFFFFFFFFFFFFC00000000000000007FFFFFFFFFFFFFFFF8000000000),
    .INIT_1B(256'h003FFFFFFFFFFFFFFFC0000000000000001FFFFFFFFFFFFFFFF8000000000000),
    .INIT_1C(256'h000FFFFFFFFFFFFFFFE0000000000000003FFFFFFFFFFFFFFFC0000000000000),
    .INIT_1D(256'h000003FFFFFFFFFFFFFFE000000000000000FFFFFFFFFFFFFFFC000000000000),
    .INIT_1E(256'h0000000007FFFFFFFFFFFFFF8000000000000007FFFFFFFFFFFFFF8000000000),
    .INIT_1F(256'h800000000000001FFFFFFFFFFFFFF800000000000001FFFFFFFFFFFFFFC00000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_049152_003 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n4242,open_n4243,open_n4244,open_n4245,open_n4246,open_n4247,open_n4248,1'b0,open_n4249}),
    .rsta(rsta),
    .doa({open_n4264,open_n4265,open_n4266,open_n4267,open_n4268,open_n4269,open_n4270,open_n4271,inst_doa_i6_003}));
  // address_offset=49152;data_offset=4;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'h000000000000000000000000000000000000000000000000000000FFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFF000000000000000000000000000000000000000000000000000),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'h00000000000000000000000000000000000000000000000000001FFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000),
    .INIT_0C(256'h000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000),
    .INIT_0E(256'h00000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000),
    .INIT_10(256'h8000000000000000000000000000000000000000000000000001FFFFFFFFFFFF),
    .INIT_11(256'h000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000000),
    .INIT_13(256'hFFFFFF000000000000000000000000000000000000000000007FFFFFFFFFFFFF),
    .INIT_14(256'h0000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'h0000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000003FFFF),
    .INIT_18(256'hFFFFFFFFFFFFF8000000000000000000000000000000000007FFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFF80000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFE0000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFC00000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFF00000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFC000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFF8000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFE00000000000000000000000000001FFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_049152_004 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n4300,open_n4301,open_n4302,open_n4303,open_n4304,open_n4305,open_n4306,1'b0,open_n4307}),
    .rsta(rsta),
    .doa({open_n4322,open_n4323,open_n4324,open_n4325,open_n4326,open_n4327,open_n4328,open_n4329,inst_doa_i6_004}));
  // address_offset=49152;data_offset=5;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'h00000000000000000000000000000000000000000000000000001FFFFFFFFFFF),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000000000),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'h00000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000),
    .INIT_11(256'h000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000),
    .INIT_14(256'h0000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFF8000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'h000000000000000000000000000000000000000000000000000000000003FFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000),
    .INIT_19(256'h000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000000000000000000),
    .INIT_1B(256'h00000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000),
    .INIT_1D(256'h000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000),
    .INIT_1F(256'h00000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_049152_005 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n4358,open_n4359,open_n4360,open_n4361,open_n4362,open_n4363,open_n4364,1'b0,open_n4365}),
    .rsta(rsta),
    .doa({open_n4380,open_n4381,open_n4382,open_n4383,open_n4384,open_n4385,open_n4386,open_n4387,inst_doa_i6_005}));
  // address_offset=49152;data_offset=6;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'h00000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'hFFFFFFFFFFFFFFF0000000000000000000000000000000000000000000000000),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'h0000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'h000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_049152_006 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n4416,open_n4417,open_n4418,open_n4419,open_n4420,open_n4421,open_n4422,1'b0,open_n4423}),
    .rsta(rsta),
    .doa({open_n4438,open_n4439,open_n4440,open_n4441,open_n4442,open_n4443,open_n4444,open_n4445,inst_doa_i6_006}));
  // address_offset=49152;data_offset=7;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000000000),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'h0000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'h000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_049152_007 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n4474,open_n4475,open_n4476,open_n4477,open_n4478,open_n4479,open_n4480,1'b0,open_n4481}),
    .rsta(rsta),
    .doa({open_n4496,open_n4497,open_n4498,open_n4499,open_n4500,open_n4501,open_n4502,open_n4503,inst_doa_i6_007}));
  // address_offset=49152;data_offset=8;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'h000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_049152_008 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n4532,open_n4533,open_n4534,open_n4535,open_n4536,open_n4537,open_n4538,1'b0,open_n4539}),
    .rsta(rsta),
    .doa({open_n4554,open_n4555,open_n4556,open_n4557,open_n4558,open_n4559,open_n4560,open_n4561,inst_doa_i6_008}));
  // address_offset=49152;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_049152_009 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n4590,open_n4591,open_n4592,open_n4593,open_n4594,open_n4595,open_n4596,1'b0,open_n4597}),
    .rsta(rsta),
    .doa({open_n4612,open_n4613,open_n4614,open_n4615,open_n4616,open_n4617,open_n4618,open_n4619,inst_doa_i6_009}));
  // address_offset=49152;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_049152_010 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n4648,open_n4649,open_n4650,open_n4651,open_n4652,open_n4653,open_n4654,1'b0,open_n4655}),
    .rsta(rsta),
    .doa({open_n4670,open_n4671,open_n4672,open_n4673,open_n4674,open_n4675,open_n4676,open_n4677,inst_doa_i6_010}));
  // address_offset=57344;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h7F01FC07F01FC07F01FC07F80FE03F80FE03F807F01FC07F01FE03F80FE01FC0),
    .INIT_01(256'h03F80FE03F80FE07F01FC07F01FC07F01FC07F01FC07F01FC07F01FC07F01FC0),
    .INIT_02(256'h0FC07F01F80FE03F01FC07F03F80FE07F01FC07F03F80FE03F81FC07F01FC07E),
    .INIT_03(256'h01F80FC07F03F81FC07E03F81FC07E03F81FC07E03F81FC07E03F81FC07F03F8),
    .INIT_04(256'h3F03F81FC0FE07F03F81FC0FE07F03F81FC0FE03F01F80FC07E03F81FC0FE07F),
    .INIT_05(256'h7F03F01F80FC0FE07E03F01F81FC0FC07E03F01F81FC0FE07E03F01F80FC07E0),
    .INIT_06(256'h03F03F81F81FC0FC0FE07E07F03F01F81F80FC0FE07E03F03F01F81FC0FC07E0),
    .INIT_07(256'h3F81F81F81F81FC0FC0FC0FE07E07E07F03F03F01F81F81FC0FC0FC07E07E07F),
    .INIT_08(256'h1F81F81F81F81F81FC0FC0FC0FC0FC0FC0FC0FE07E07E07E07E07F03F03F03F0),
    .INIT_09(256'hC0FC0FC1F81F81F81F81F81F81F81F81F81F81F81F81F81F81F81F81F81F81F8),
    .INIT_0A(256'h0FC0FC0F81F81F81F81F03F03F03F03F07E07E07E07E07E07C0FC0FC0FC0FC0F),
    .INIT_0B(256'h0FC0FC1F81F83F03F03E07E07E0FC0FC0FC1F81F81F03F03F03F07E07E07E0FC),
    .INIT_0C(256'hC0F81F83F03F07E07C0FC0F81F81F03F03E07E0FC0FC1F81F81F03F03E07E07C),
    .INIT_0D(256'h1F03F07E07C0FC1F81F03E07E0FC0F81F83F03E07E07C0FC1F81F03F07E07C0F),
    .INIT_0E(256'h7E0FC1F83F03E07C0FC1F83F03E07C0FC1F83F03E07C0FC1F83F03E07E0FC0F8),
    .INIT_0F(256'h3F07E0FC1F83F07E0FC1F83F07E07C0F81F03E07C0FC1F83F07E0FC0F81F03E0),
    .INIT_10(256'h03E07C1F83F07E0FC1F83F07E0FC1F83E07C0F81F03E07C0F81F03E07C0F81F0),
    .INIT_11(256'h7C0F83F07E0F81F03E07C1F83F07E0F81F03E07C1F83F07E0FC1F03E07C0F81F),
    .INIT_12(256'hE07C0F83F07C0F81F07E0F81F03E0FC1F03E07C1F83F07C0F81F07E0FC1F03E0),
    .INIT_13(256'hE0FC1F03E0FC1F03E0FC1F03E0FC1F03E0FC1F03E0FC1F03E0FC1F83E07C1F83),
    .INIT_14(256'hF03E0F81F07E0F83F07C0F83F07C1F83E07C1F83E07C1F03E0FC1F03E0FC1F03),
    .INIT_15(256'h3E07C1F03E0F81F07C0F83E07C1F83E0FC1F07E0F81F07C0F83E07C1F83E0FC1),
    .INIT_16(256'hC1F07C0F83E07C1F07E0F83F07C1F83E0F81F07C0F83E07C1F03E0F81F07C0F8),
    .INIT_17(256'h3F07C1F03E0F83F07C1F03E0F83F07C1F03E0F83F07C1F03E0F81F07C1F83E0F),
    .INIT_18(256'hF03E0F83E07C1F07E0F83E0FC1F07C1F83E0F81F07C1F83E0F83F07C1F03E0F8),
    .INIT_19(256'hC0F83E0F83F07C1F07E0F83E0FC1F07C1F03E0F83E07C1F07C0F83E0F81F07C1),
    .INIT_1A(256'h81F07C1F07C0F83E0F83F07C1F07C0F83E0F83F07C1F07C0F83E0F83F07C1F07),
    .INIT_1B(256'h83E0FC1F07C1F07E0F83E0F83F07C1F07C1F83E0F83E0FC1F07C1F07E0F83E0F),
    .INIT_1C(256'h81F07C1F07C1F83E0F83E0F81F07C1F07C1F83E0F83E0F81F07C1F07C1F83E0F),
    .INIT_1D(256'hC1F03E0F83E0F83E07C1F07C1F07C0F83E0F83E0FC1F07C1F07C1F83E0F83E0F),
    .INIT_1E(256'hE0FC1F07C1F07C1F03E0F83E0F83E07C1F07C1F07C0F83E0F83E0F81F07C1F07),
    .INIT_1F(256'hF83E0F83E0F83F07C1F07C1F07C0F83E0F83E0F81F07C1F07C1F07E0F83E0F83),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_057344_000 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n4706,open_n4707,open_n4708,open_n4709,open_n4710,open_n4711,open_n4712,1'b0,open_n4713}),
    .rsta(rsta),
    .doa({open_n4728,open_n4729,open_n4730,open_n4731,open_n4732,open_n4733,open_n4734,open_n4735,inst_doa_i7_000}));
  // address_offset=57344;data_offset=1;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h7FFE0007FFE0007FFE0007FFF0003FFF0003FFF8001FFF8001FFFC000FFFE000),
    .INIT_01(256'h03FFF0003FFF0007FFE0007FFE0007FFE0007FFE0007FFE0007FFE0007FFE000),
    .INIT_02(256'hF0007FFE000FFFC001FFF8003FFF0007FFE0007FFC000FFFC001FFF8001FFF80),
    .INIT_03(256'h01FFF0007FFC001FFF8003FFE0007FFC001FFF8003FFE0007FFC001FFF8003FF),
    .INIT_04(256'h3FFC001FFF0007FFC001FFF0007FFC001FFF0003FFE000FFF8003FFE000FFF80),
    .INIT_05(256'h7FFC001FFF000FFF8003FFE001FFF0007FFC001FFE000FFF8003FFE000FFF800),
    .INIT_06(256'h03FFC001FFE000FFF0007FF8003FFE001FFF000FFF8003FFC001FFE000FFF800),
    .INIT_07(256'hC001FFE001FFE000FFF000FFF8007FF8003FFC001FFE001FFF000FFF8007FF80),
    .INIT_08(256'h1FFE001FFE001FFE000FFF000FFF000FFF000FFF8007FF8007FF8003FFC003FF),
    .INIT_09(256'hFF000FFE001FFE001FFE001FFE001FFE001FFE001FFE001FFE001FFE001FFE00),
    .INIT_0A(256'hF000FFF001FFE001FFE003FFC003FFC007FF8007FF8007FF800FFF000FFF000F),
    .INIT_0B(256'hF000FFE001FFC003FFC007FF800FFF000FFE001FFE003FFC003FF8007FF800FF),
    .INIT_0C(256'hFF001FFC003FF8007FF000FFE001FFC003FF800FFF001FFE001FFC003FF8007F),
    .INIT_0D(256'h1FFC007FF800FFE001FFC007FF000FFE003FFC007FF800FFE001FFC007FF800F),
    .INIT_0E(256'h800FFE003FFC007FF001FFC003FF800FFE003FFC007FF001FFC003FF800FFF00),
    .INIT_0F(256'h3FF800FFE003FF800FFE003FF8007FF001FFC007FF001FFC007FF000FFE003FF),
    .INIT_10(256'hFC007FE003FF800FFE003FF800FFE003FF800FFE003FF800FFE003FF800FFE00),
    .INIT_11(256'h800FFC007FF001FFC007FE003FF800FFE003FF801FFC007FF001FFC007FF001F),
    .INIT_12(256'h007FF003FF800FFE007FF001FFC00FFE003FF801FFC007FF001FF800FFE003FF),
    .INIT_13(256'h00FFE003FF001FFC00FFE003FF001FFC00FFE003FF001FFC00FFE003FF801FFC),
    .INIT_14(256'h003FF001FF800FFC007FF003FF801FFC007FE003FF801FFC00FFE003FF001FFC),
    .INIT_15(256'hC007FE003FF001FF800FFC007FE003FF001FF800FFE007FF003FF801FFC00FFE),
    .INIT_16(256'hFE007FF003FF801FF800FFC007FE003FF001FF800FFC007FE003FF001FF800FF),
    .INIT_17(256'h3FF801FFC00FFC007FE003FF003FF801FFC00FFC007FE003FF001FF801FFC00F),
    .INIT_18(256'h003FF003FF801FF800FFC00FFE007FE003FF001FF801FFC00FFC007FE003FF00),
    .INIT_19(256'hFF003FF003FF801FF800FFC00FFE007FE003FF003FF801FF800FFC00FFE007FE),
    .INIT_1A(256'h01FF801FF800FFC00FFC007FE007FF003FF003FF801FF800FFC00FFC007FE007),
    .INIT_1B(256'hFC00FFE007FE007FF003FF003FF801FF801FFC00FFC00FFE007FE007FF003FF0),
    .INIT_1C(256'h01FF801FF801FFC00FFC00FFE007FE007FE003FF003FF001FF801FF801FFC00F),
    .INIT_1D(256'hFE003FF003FF003FF801FF801FF800FFC00FFC00FFE007FE007FE003FF003FF0),
    .INIT_1E(256'h00FFE007FE007FE003FF003FF003FF801FF801FF800FFC00FFC00FFE007FE007),
    .INIT_1F(256'hFFC00FFC00FFC007FE007FE007FF003FF003FF001FF801FF801FF800FFC00FFC),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_057344_001 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n4764,open_n4765,open_n4766,open_n4767,open_n4768,open_n4769,open_n4770,1'b0,open_n4771}),
    .rsta(rsta),
    .doa({open_n4786,open_n4787,open_n4788,open_n4789,open_n4790,open_n4791,open_n4792,open_n4793,inst_doa_i7_001}));
  // address_offset=57344;data_offset=2;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h80000007FFFFFF80000007FFFFFFC0000003FFFFFFE0000001FFFFFFF0000000),
    .INIT_01(256'h03FFFFFFC0000007FFFFFF80000007FFFFFF80000007FFFFFF80000007FFFFFF),
    .INIT_02(256'hFFFF8000000FFFFFFE0000003FFFFFF80000007FFFFFF0000001FFFFFFE00000),
    .INIT_03(256'hFE0000007FFFFFE0000003FFFFFF8000001FFFFFFC0000007FFFFFE0000003FF),
    .INIT_04(256'hC000001FFFFFF8000001FFFFFF8000001FFFFFFC000000FFFFFFC000000FFFFF),
    .INIT_05(256'h8000001FFFFFF0000003FFFFFE0000007FFFFFE000000FFFFFFC000000FFFFFF),
    .INIT_06(256'hFC000001FFFFFF0000007FFFFFC000001FFFFFF0000003FFFFFE000000FFFFFF),
    .INIT_07(256'hFFFE000001FFFFFF000000FFFFFF8000003FFFFFE000001FFFFFF0000007FFFF),
    .INIT_08(256'h1FFFFFE000001FFFFFF000000FFFFFF000000FFFFFF8000007FFFFFC000003FF),
    .INIT_09(256'h00000FFFFFE000001FFFFFE000001FFFFFE000001FFFFFE000001FFFFFE00000),
    .INIT_0A(256'hFFFF000001FFFFFE000003FFFFFC000007FFFFF8000007FFFFF000000FFFFFF0),
    .INIT_0B(256'h0000FFFFFE000003FFFFF800000FFFFFF000001FFFFFC000003FFFFF800000FF),
    .INIT_0C(256'hFFFFE000003FFFFF800000FFFFFE000003FFFFF000001FFFFFE000003FFFFF80),
    .INIT_0D(256'hE000007FFFFF000001FFFFF800000FFFFFC000007FFFFF000001FFFFF800000F),
    .INIT_0E(256'h000FFFFFC000007FFFFE000003FFFFF000003FFFFF800001FFFFFC00000FFFFF),
    .INIT_0F(256'h3FFFFF000003FFFFF000003FFFFF800001FFFFF800001FFFFF800000FFFFFC00),
    .INIT_10(256'hFFFF800003FFFFF000003FFFFF000003FFFFF000003FFFFF000003FFFFF00000),
    .INIT_11(256'hFFF000007FFFFE000007FFFFC00000FFFFFC00001FFFFF800001FFFFF800001F),
    .INIT_12(256'hFF800003FFFFF000007FFFFE00000FFFFFC00001FFFFF800001FFFFF000003FF),
    .INIT_13(256'hFF000003FFFFE00000FFFFFC00001FFFFF000003FFFFE00000FFFFFC00001FFF),
    .INIT_14(256'hFFC00001FFFFF000007FFFFC00001FFFFF800003FFFFE00000FFFFFC00001FFF),
    .INIT_15(256'hFFF800003FFFFE00000FFFFF800003FFFFE00000FFFFF800003FFFFE00000FFF),
    .INIT_16(256'hFFFF800003FFFFE00000FFFFF800003FFFFE00000FFFFF800003FFFFE00000FF),
    .INIT_17(256'h3FFFFE00000FFFFF800003FFFFC00001FFFFF000007FFFFC00001FFFFE00000F),
    .INIT_18(256'h003FFFFC00001FFFFF00000FFFFF800003FFFFE00001FFFFF000007FFFFC0000),
    .INIT_19(256'h00003FFFFC00001FFFFF00000FFFFF800003FFFFC00001FFFFF00000FFFFF800),
    .INIT_1A(256'hFE00001FFFFF00000FFFFF800007FFFFC00003FFFFE00000FFFFF000007FFFF8),
    .INIT_1B(256'hFFFF000007FFFF800003FFFFC00001FFFFE00000FFFFF000007FFFF800003FFF),
    .INIT_1C(256'h01FFFFE00001FFFFF00000FFFFF800007FFFFC00003FFFFE00001FFFFE00000F),
    .INIT_1D(256'h00003FFFFC00003FFFFE00001FFFFF00000FFFFF000007FFFF800003FFFFC000),
    .INIT_1E(256'hFF000007FFFF800003FFFFC00003FFFFE00001FFFFF00000FFFFF000007FFFF8),
    .INIT_1F(256'hFFFFF00000FFFFF800007FFFF800003FFFFC00001FFFFE00001FFFFF00000FFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_057344_002 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n4822,open_n4823,open_n4824,open_n4825,open_n4826,open_n4827,open_n4828,1'b0,open_n4829}),
    .rsta(rsta),
    .doa({open_n4844,open_n4845,open_n4846,open_n4847,open_n4848,open_n4849,open_n4850,open_n4851,inst_doa_i7_002}));
  // address_offset=57344;data_offset=3;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFF800000000000007FFFFFFFFFFFFFC00000000000001FFFFFFFFFFFFFF),
    .INIT_01(256'h03FFFFFFFFFFFFF800000000000007FFFFFFFFFFFFF800000000000007FFFFFF),
    .INIT_02(256'h00000000000FFFFFFFFFFFFFC00000000000007FFFFFFFFFFFFE000000000000),
    .INIT_03(256'hFFFFFFFF80000000000003FFFFFFFFFFFFE00000000000007FFFFFFFFFFFFC00),
    .INIT_04(256'h0000001FFFFFFFFFFFFE0000000000001FFFFFFFFFFFFF0000000000000FFFFF),
    .INIT_05(256'hFFFFFFE0000000000003FFFFFFFFFFFF8000000000000FFFFFFFFFFFFF000000),
    .INIT_06(256'h00000001FFFFFFFFFFFF8000000000001FFFFFFFFFFFFC000000000000FFFFFF),
    .INIT_07(256'hFFFFFFFFFE000000000000FFFFFFFFFFFFC000000000001FFFFFFFFFFFF80000),
    .INIT_08(256'hE000000000001FFFFFFFFFFFF000000000000FFFFFFFFFFFF8000000000003FF),
    .INIT_09(256'h00000FFFFFFFFFFFE000000000001FFFFFFFFFFFE000000000001FFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFE000000000003FFFFFFFFFFF8000000000007FFFFFFFFFFF0000000),
    .INIT_0B(256'hFFFF000000000003FFFFFFFFFFF000000000001FFFFFFFFFFFC00000000000FF),
    .INIT_0C(256'h00000000003FFFFFFFFFFF000000000003FFFFFFFFFFE000000000003FFFFFFF),
    .INIT_0D(256'h0000007FFFFFFFFFFE00000000000FFFFFFFFFFF800000000001FFFFFFFFFFF0),
    .INIT_0E(256'h000FFFFFFFFFFF800000000003FFFFFFFFFFC00000000001FFFFFFFFFFF00000),
    .INIT_0F(256'h3FFFFFFFFFFC00000000003FFFFFFFFFFE00000000001FFFFFFFFFFF00000000),
    .INIT_10(256'hFFFFFFFFFC00000000003FFFFFFFFFFC00000000003FFFFFFFFFFC0000000000),
    .INIT_11(256'hFFFFFFFF800000000007FFFFFFFFFF00000000001FFFFFFFFFFE00000000001F),
    .INIT_12(256'hFFFFFFFC00000000007FFFFFFFFFF00000000001FFFFFFFFFFE00000000003FF),
    .INIT_13(256'hFFFFFFFC0000000000FFFFFFFFFFE00000000003FFFFFFFFFF00000000001FFF),
    .INIT_14(256'hFFFFFFFE00000000007FFFFFFFFFE00000000003FFFFFFFFFF00000000001FFF),
    .INIT_15(256'hFFFFFFFFC0000000000FFFFFFFFFFC0000000000FFFFFFFFFFC0000000000FFF),
    .INIT_16(256'hFFFFFFFFFC0000000000FFFFFFFFFFC0000000000FFFFFFFFFFC0000000000FF),
    .INIT_17(256'h3FFFFFFFFFF00000000003FFFFFFFFFE00000000007FFFFFFFFFE0000000000F),
    .INIT_18(256'h003FFFFFFFFFE0000000000FFFFFFFFFFC0000000001FFFFFFFFFF8000000000),
    .INIT_19(256'h00003FFFFFFFFFE0000000000FFFFFFFFFFC0000000001FFFFFFFFFF00000000),
    .INIT_1A(256'h0000001FFFFFFFFFF00000000007FFFFFFFFFC0000000000FFFFFFFFFF800000),
    .INIT_1B(256'h0000000007FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFFFFFFC000),
    .INIT_1C(256'hFE0000000001FFFFFFFFFF00000000007FFFFFFFFFC0000000001FFFFFFFFFF0),
    .INIT_1D(256'hFFFFC0000000003FFFFFFFFFE0000000000FFFFFFFFFF80000000003FFFFFFFF),
    .INIT_1E(256'hFFFFFFF80000000003FFFFFFFFFC0000000001FFFFFFFFFF00000000007FFFFF),
    .INIT_1F(256'hFFFFFFFFFF00000000007FFFFFFFFFC0000000001FFFFFFFFFE0000000000FFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_057344_003 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n4880,open_n4881,open_n4882,open_n4883,open_n4884,open_n4885,open_n4886,1'b0,open_n4887}),
    .rsta(rsta),
    .doa({open_n4902,open_n4903,open_n4904,open_n4905,open_n4906,open_n4907,open_n4908,open_n4909,inst_doa_i7_003}));
  // address_offset=57344;data_offset=4;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000001FFFFFFFFFFFFFF),
    .INIT_01(256'h03FFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000007FFFFFF),
    .INIT_02(256'h00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000000000000000),
    .INIT_03(256'h0000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000),
    .INIT_04(256'hFFFFFFE00000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFF00000),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFC0000000000000000000000000FFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'h00000001FFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000FFFFFF),
    .INIT_07(256'h0000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000),
    .INIT_08(256'hFFFFFFFFFFFFE000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFC00),
    .INIT_09(256'h00000FFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000001FFFFFFFFFFF),
    .INIT_0A(256'h0000000000000000000003FFFFFFFFFFFFFFFFFFFFFFF8000000000000000000),
    .INIT_0B(256'hFFFFFFFFFFFFFFFC00000000000000000000001FFFFFFFFFFFFFFFFFFFFFFF00),
    .INIT_0C(256'h00000000003FFFFFFFFFFFFFFFFFFFFFFC00000000000000000000003FFFFFFF),
    .INIT_0D(256'hFFFFFF80000000000000000000000FFFFFFFFFFFFFFFFFFFFFFE000000000000),
    .INIT_0E(256'h000FFFFFFFFFFFFFFFFFFFFFFC0000000000000000000001FFFFFFFFFFFFFFFF),
    .INIT_0F(256'hC0000000000000000000003FFFFFFFFFFFFFFFFFFFFFE0000000000000000000),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFC0000000000000000000003FFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h00000000000000000007FFFFFFFFFFFFFFFFFFFFE0000000000000000000001F),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFF8000000000000000000001FFFFFFFFFFFFFFFFFFFFFC00),
    .INIT_13(256'h000000000000000000FFFFFFFFFFFFFFFFFFFFFC000000000000000000001FFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFF8000000000000000000003FFFFFFFFFFFFFFFFFFFFE000),
    .INIT_15(256'h0000000000000000000FFFFFFFFFFFFFFFFFFFFF000000000000000000000FFF),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFF000000000000000000000FFFFFFFFFFFFFFFFFFFFF00),
    .INIT_17(256'hC000000000000000000003FFFFFFFFFFFFFFFFFFFF800000000000000000000F),
    .INIT_18(256'h003FFFFFFFFFFFFFFFFFFFF000000000000000000001FFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFFE000000000000000000),
    .INIT_1A(256'h0000001FFFFFFFFFFFFFFFFFFFF800000000000000000000FFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFF800000000000000000001FFFFFFFFFFFFFFFFFFFF80000000000000),
    .INIT_1C(256'h000000000001FFFFFFFFFFFFFFFFFFFF800000000000000000001FFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFC00000000000000000000FFFFFFFFFFFFFFFFFFFFC00000000),
    .INIT_1E(256'h000000000000000003FFFFFFFFFFFFFFFFFFFE000000000000000000007FFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFF800000000000000000001FFFFFFFFFFFFFFFFFFFF000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_057344_004 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n4938,open_n4939,open_n4940,open_n4941,open_n4942,open_n4943,open_n4944,1'b0,open_n4945}),
    .rsta(rsta),
    .doa({open_n4960,open_n4961,open_n4962,open_n4963,open_n4964,open_n4965,open_n4966,open_n4967,inst_doa_i7_004}));
  // address_offset=57344;data_offset=5;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000),
    .INIT_01(256'hFC00000000000000000000000000000000000000000000000000000007FFFFFF),
    .INIT_02(256'h00000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000),
    .INIT_04(256'h000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000),
    .INIT_06(256'hFFFFFFFE00000000000000000000000000000000000000000000000000FFFFFF),
    .INIT_07(256'h0000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000),
    .INIT_09(256'hFFFFF000000000000000000000000000000000000000000000001FFFFFFFFFFF),
    .INIT_0A(256'h0000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000),
    .INIT_0C(256'hFFFFFFFFFFC0000000000000000000000000000000000000000000003FFFFFFF),
    .INIT_0D(256'h00000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'h000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h00000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFF0000000000000000000000000000000000000000001FFF),
    .INIT_14(256'h0000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'h0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFC00000000000000000000000000000000000000000F),
    .INIT_18(256'hFFC00000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'h0000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'h0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000000),
    .INIT_1C(256'hFFFFFFFFFFFE00000000000000000000000000000000000000001FFFFFFFFFFF),
    .INIT_1D(256'h00000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'h000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_057344_005 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n4996,open_n4997,open_n4998,open_n4999,open_n5000,open_n5001,open_n5002,1'b0,open_n5003}),
    .rsta(rsta),
    .doa({open_n5018,open_n5019,open_n5020,open_n5021,open_n5022,open_n5023,open_n5024,open_n5025,inst_doa_i7_005}));
  // address_offset=57344;data_offset=6;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000007FFFFFF),
    .INIT_02(256'hFFFFFFFFFFF00000000000000000000000000000000000000000000000000000),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'h000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000),
    .INIT_07(256'h0000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000),
    .INIT_0A(256'h0000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000),
    .INIT_0D(256'h00000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFF0000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'h0000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFF800000000000000000000000000000000000000000000),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000001FFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000),
    .INIT_15(256'h0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0),
    .INIT_18(256'h00000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000),
    .INIT_1A(256'h0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000),
    .INIT_1D(256'h00000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFC0000000000000000000000000000000000000000000000),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_057344_006 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n5054,open_n5055,open_n5056,open_n5057,open_n5058,open_n5059,open_n5060,1'b0,open_n5061}),
    .rsta(rsta),
    .doa({open_n5076,open_n5077,open_n5078,open_n5079,open_n5080,open_n5081,open_n5082,open_n5083,inst_doa_i7_006}));
  // address_offset=57344;data_offset=7;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'h000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'h0000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000000),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'h0000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'h0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000000000),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'h0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_057344_007 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n5112,open_n5113,open_n5114,open_n5115,open_n5116,open_n5117,open_n5118,1'b0,open_n5119}),
    .rsta(rsta),
    .doa({open_n5134,open_n5135,open_n5136,open_n5137,open_n5138,open_n5139,open_n5140,open_n5141,inst_doa_i7_007}));
  // address_offset=57344;data_offset=8;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'h0000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'h0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'hFFFFFFE000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_057344_008 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n5170,open_n5171,open_n5172,open_n5173,open_n5174,open_n5175,open_n5176,1'b0,open_n5177}),
    .rsta(rsta),
    .doa({open_n5192,open_n5193,open_n5194,open_n5195,open_n5196,open_n5197,open_n5198,open_n5199,inst_doa_i7_008}));
  // address_offset=57344;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'h0000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_057344_009 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n5228,open_n5229,open_n5230,open_n5231,open_n5232,open_n5233,open_n5234,1'b0,open_n5235}),
    .rsta(rsta),
    .doa({open_n5250,open_n5251,open_n5252,open_n5253,open_n5254,open_n5255,open_n5256,open_n5257,inst_doa_i7_009}));
  // address_offset=57344;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_057344_010 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n5286,open_n5287,open_n5288,open_n5289,open_n5290,open_n5291,open_n5292,1'b0,open_n5293}),
    .rsta(rsta),
    .doa({open_n5308,open_n5309,open_n5310,open_n5311,open_n5312,open_n5313,open_n5314,open_n5315,inst_doa_i7_010}));
  // address_offset=57344;data_offset=11;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_057344_011 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n5344,open_n5345,open_n5346,open_n5347,open_n5348,open_n5349,open_n5350,1'b0,open_n5351}),
    .rsta(rsta),
    .doa({open_n5366,open_n5367,open_n5368,open_n5369,open_n5370,open_n5371,open_n5372,open_n5373,inst_doa_i7_011}));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_0  (
    .i0(inst_doa_i0_000),
    .i1(inst_doa_i1_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_0 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_1  (
    .i0(inst_doa_i2_000),
    .i1(inst_doa_i3_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_1 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_2  (
    .i0(inst_doa_i4_000),
    .i1(inst_doa_i5_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_2 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_3  (
    .i0(inst_doa_i6_000),
    .i1(inst_doa_i7_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_3 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b0/B0_0 ),
    .i1(\inst_doa_mux_b0/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_0 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b0/B0_2 ),
    .i1(\inst_doa_mux_b0/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_1 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b0/B1_0 ),
    .i1(\inst_doa_mux_b0/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[0]));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_0  (
    .i0(inst_doa_i0_001),
    .i1(inst_doa_i1_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_0 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_1  (
    .i0(inst_doa_i2_001),
    .i1(inst_doa_i3_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_1 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_2  (
    .i0(inst_doa_i4_001),
    .i1(inst_doa_i5_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_2 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_3  (
    .i0(inst_doa_i6_001),
    .i1(inst_doa_i7_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_3 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b1/B0_0 ),
    .i1(\inst_doa_mux_b1/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_0 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b1/B0_2 ),
    .i1(\inst_doa_mux_b1/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_1 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b1/B1_0 ),
    .i1(\inst_doa_mux_b1/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[1]));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_0_0  (
    .i0(inst_doa_i0_010),
    .i1(inst_doa_i1_010),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b10/B0_0 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_0_1  (
    .i0(inst_doa_i2_010),
    .i1(inst_doa_i3_010),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b10/B0_1 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_0_2  (
    .i0(inst_doa_i4_010),
    .i1(inst_doa_i5_010),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b10/B0_2 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_0_3  (
    .i0(inst_doa_i6_010),
    .i1(inst_doa_i7_010),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b10/B0_3 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b10/B0_0 ),
    .i1(\inst_doa_mux_b10/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b10/B1_0 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b10/B0_2 ),
    .i1(\inst_doa_mux_b10/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b10/B1_1 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b10/B1_0 ),
    .i1(\inst_doa_mux_b10/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[10]));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_0_0  (
    .i0(inst_doa_i0_011),
    .i1(inst_doa_i1_010),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b11/B0_0 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_0_1  (
    .i0(inst_doa_i2_010),
    .i1(inst_doa_i3_011),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b11/B0_1 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_0_2  (
    .i0(inst_doa_i4_011),
    .i1(inst_doa_i5_010),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b11/B0_2 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_0_3  (
    .i0(inst_doa_i6_010),
    .i1(inst_doa_i7_011),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b11/B0_3 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b11/B0_0 ),
    .i1(\inst_doa_mux_b11/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b11/B1_0 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b11/B0_2 ),
    .i1(\inst_doa_mux_b11/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b11/B1_1 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b11/B1_0 ),
    .i1(\inst_doa_mux_b11/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[11]));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_0  (
    .i0(inst_doa_i0_002),
    .i1(inst_doa_i1_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_0 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_1  (
    .i0(inst_doa_i2_002),
    .i1(inst_doa_i3_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_1 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_2  (
    .i0(inst_doa_i4_002),
    .i1(inst_doa_i5_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_2 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_3  (
    .i0(inst_doa_i6_002),
    .i1(inst_doa_i7_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_3 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b2/B0_0 ),
    .i1(\inst_doa_mux_b2/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_0 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b2/B0_2 ),
    .i1(\inst_doa_mux_b2/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_1 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b2/B1_0 ),
    .i1(\inst_doa_mux_b2/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[2]));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_0  (
    .i0(inst_doa_i0_003),
    .i1(inst_doa_i1_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_0 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_1  (
    .i0(inst_doa_i2_003),
    .i1(inst_doa_i3_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_1 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_2  (
    .i0(inst_doa_i4_003),
    .i1(inst_doa_i5_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_2 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_3  (
    .i0(inst_doa_i6_003),
    .i1(inst_doa_i7_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_3 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b3/B0_0 ),
    .i1(\inst_doa_mux_b3/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_0 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b3/B0_2 ),
    .i1(\inst_doa_mux_b3/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_1 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b3/B1_0 ),
    .i1(\inst_doa_mux_b3/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[3]));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_0  (
    .i0(inst_doa_i0_004),
    .i1(inst_doa_i1_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_0 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_1  (
    .i0(inst_doa_i2_004),
    .i1(inst_doa_i3_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_1 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_2  (
    .i0(inst_doa_i4_004),
    .i1(inst_doa_i5_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_2 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_3  (
    .i0(inst_doa_i6_004),
    .i1(inst_doa_i7_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_3 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b4/B0_0 ),
    .i1(\inst_doa_mux_b4/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_0 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b4/B0_2 ),
    .i1(\inst_doa_mux_b4/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_1 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b4/B1_0 ),
    .i1(\inst_doa_mux_b4/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[4]));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_0  (
    .i0(inst_doa_i0_005),
    .i1(inst_doa_i1_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_0 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_1  (
    .i0(inst_doa_i2_005),
    .i1(inst_doa_i3_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_1 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_2  (
    .i0(inst_doa_i4_005),
    .i1(inst_doa_i5_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_2 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_3  (
    .i0(inst_doa_i6_005),
    .i1(inst_doa_i7_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_3 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b5/B0_0 ),
    .i1(\inst_doa_mux_b5/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_0 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b5/B0_2 ),
    .i1(\inst_doa_mux_b5/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_1 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b5/B1_0 ),
    .i1(\inst_doa_mux_b5/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[5]));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_0  (
    .i0(inst_doa_i0_006),
    .i1(inst_doa_i1_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_0 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_1  (
    .i0(inst_doa_i2_006),
    .i1(inst_doa_i3_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_1 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_2  (
    .i0(inst_doa_i4_006),
    .i1(inst_doa_i5_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_2 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_3  (
    .i0(inst_doa_i6_006),
    .i1(inst_doa_i7_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_3 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b6/B0_0 ),
    .i1(\inst_doa_mux_b6/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_0 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b6/B0_2 ),
    .i1(\inst_doa_mux_b6/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_1 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b6/B1_0 ),
    .i1(\inst_doa_mux_b6/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[6]));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_0  (
    .i0(inst_doa_i0_007),
    .i1(inst_doa_i1_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_0 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_1  (
    .i0(inst_doa_i2_007),
    .i1(inst_doa_i3_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_1 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_2  (
    .i0(inst_doa_i4_007),
    .i1(inst_doa_i5_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_2 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_3  (
    .i0(inst_doa_i6_007),
    .i1(inst_doa_i7_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_3 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b7/B0_0 ),
    .i1(\inst_doa_mux_b7/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_0 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b7/B0_2 ),
    .i1(\inst_doa_mux_b7/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_1 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b7/B1_0 ),
    .i1(\inst_doa_mux_b7/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[7]));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_0  (
    .i0(inst_doa_i0_008),
    .i1(inst_doa_i1_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_0 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_1  (
    .i0(inst_doa_i2_008),
    .i1(inst_doa_i3_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_1 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_2  (
    .i0(inst_doa_i4_008),
    .i1(inst_doa_i5_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_2 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_3  (
    .i0(inst_doa_i6_008),
    .i1(inst_doa_i7_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_3 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b8/B0_0 ),
    .i1(\inst_doa_mux_b8/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_0 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b8/B0_2 ),
    .i1(\inst_doa_mux_b8/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_1 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b8/B1_0 ),
    .i1(\inst_doa_mux_b8/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[8]));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_0_0  (
    .i0(inst_doa_i0_009),
    .i1(inst_doa_i1_009),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b9/B0_0 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_0_1  (
    .i0(inst_doa_i2_009),
    .i1(inst_doa_i3_009),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b9/B0_1 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_0_2  (
    .i0(inst_doa_i4_009),
    .i1(inst_doa_i5_009),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b9/B0_2 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_0_3  (
    .i0(inst_doa_i6_009),
    .i1(inst_doa_i7_009),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b9/B0_3 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b9/B0_0 ),
    .i1(\inst_doa_mux_b9/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b9/B1_0 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b9/B0_2 ),
    .i1(\inst_doa_mux_b9/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b9/B1_1 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b9/B1_0 ),
    .i1(\inst_doa_mux_b9/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[9]));

endmodule 

module AL_DFF_X
  (
  ar,
  as,
  clk,
  d,
  en,
  sr,
  ss,
  q
  );

  input ar;
  input as;
  input clk;
  input d;
  input en;
  input sr;
  input ss;
  output q;

  wire enout;
  wire srout;
  wire ssout;

  AL_MUX u_en (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_MUX u_reset (
    .i0(ssout),
    .i1(1'b0),
    .sel(sr),
    .o(srout));
  AL_DFF u_seq (
    .clk(clk),
    .d(srout),
    .reset(ar),
    .set(as),
    .q(q));
  AL_MUX u_set (
    .i0(enout),
    .i1(1'b1),
    .sel(ss),
    .o(ssout));

endmodule 

module AL_MUX
  (
  input i0,
  input i1,
  input sel,
  output o
  );

  wire not_sel, sel_i0, sel_i1;
  not u0 (not_sel, sel);
  and u1 (sel_i1, sel, i1);
  and u2 (sel_i0, not_sel, i0);
  or u3 (o, sel_i1, sel_i0);

endmodule

module AL_DFF
  (
  input reset,
  input set,
  input clk,
  input d,
  output reg q
  );

  parameter INI = 1'b0;

  // synthesis translate_off
  tri0 gsrn = glbl.gsrn;

  always @(gsrn)
  begin
    if(!gsrn)
      assign q = INI;
    else
      deassign q;
  end
  // synthesis translate_on

  always @(posedge reset or posedge set or posedge clk)
  begin
    if (reset)
      q <= 1'b0;
    else if (set)
      q <= 1'b1;
    else
      q <= d;
  end

endmodule

