// Verilog netlist created by TD v5.0.30786
// Wed Aug 24 13:29:02 2022

`timescale 1ns / 1ps
module ROM_Cos_table  // ROM_Cos_table.v(14)
  (
  addra,
  clka,
  rsta,
  doa
  );

  input [15:0] addra;  // ROM_Cos_table.v(18)
  input clka;  // ROM_Cos_table.v(19)
  input rsta;  // ROM_Cos_table.v(20)
  output [11:0] doa;  // ROM_Cos_table.v(16)

  wire [0:5] addra_piped;
  wire  \inst_doa_mux_b0/B0_0 ;
  wire  \inst_doa_mux_b0/B0_1 ;
  wire  \inst_doa_mux_b0/B0_10 ;
  wire  \inst_doa_mux_b0/B0_11 ;
  wire  \inst_doa_mux_b0/B0_12 ;
  wire  \inst_doa_mux_b0/B0_13 ;
  wire  \inst_doa_mux_b0/B0_14 ;
  wire  \inst_doa_mux_b0/B0_15 ;
  wire  \inst_doa_mux_b0/B0_16 ;
  wire  \inst_doa_mux_b0/B0_17 ;
  wire  \inst_doa_mux_b0/B0_18 ;
  wire  \inst_doa_mux_b0/B0_19 ;
  wire  \inst_doa_mux_b0/B0_2 ;
  wire  \inst_doa_mux_b0/B0_20 ;
  wire  \inst_doa_mux_b0/B0_21 ;
  wire  \inst_doa_mux_b0/B0_22 ;
  wire  \inst_doa_mux_b0/B0_23 ;
  wire  \inst_doa_mux_b0/B0_24 ;
  wire  \inst_doa_mux_b0/B0_25 ;
  wire  \inst_doa_mux_b0/B0_26 ;
  wire  \inst_doa_mux_b0/B0_27 ;
  wire  \inst_doa_mux_b0/B0_28 ;
  wire  \inst_doa_mux_b0/B0_29 ;
  wire  \inst_doa_mux_b0/B0_3 ;
  wire  \inst_doa_mux_b0/B0_30 ;
  wire  \inst_doa_mux_b0/B0_31 ;
  wire  \inst_doa_mux_b0/B0_4 ;
  wire  \inst_doa_mux_b0/B0_5 ;
  wire  \inst_doa_mux_b0/B0_6 ;
  wire  \inst_doa_mux_b0/B0_7 ;
  wire  \inst_doa_mux_b0/B0_8 ;
  wire  \inst_doa_mux_b0/B0_9 ;
  wire  \inst_doa_mux_b0/B1_0 ;
  wire  \inst_doa_mux_b0/B1_1 ;
  wire  \inst_doa_mux_b0/B1_10 ;
  wire  \inst_doa_mux_b0/B1_11 ;
  wire  \inst_doa_mux_b0/B1_12 ;
  wire  \inst_doa_mux_b0/B1_13 ;
  wire  \inst_doa_mux_b0/B1_14 ;
  wire  \inst_doa_mux_b0/B1_15 ;
  wire  \inst_doa_mux_b0/B1_2 ;
  wire  \inst_doa_mux_b0/B1_3 ;
  wire  \inst_doa_mux_b0/B1_4 ;
  wire  \inst_doa_mux_b0/B1_5 ;
  wire  \inst_doa_mux_b0/B1_6 ;
  wire  \inst_doa_mux_b0/B1_7 ;
  wire  \inst_doa_mux_b0/B1_8 ;
  wire  \inst_doa_mux_b0/B1_9 ;
  wire  \inst_doa_mux_b0/B2_0 ;
  wire  \inst_doa_mux_b0/B2_1 ;
  wire  \inst_doa_mux_b0/B2_2 ;
  wire  \inst_doa_mux_b0/B2_3 ;
  wire  \inst_doa_mux_b0/B2_4 ;
  wire  \inst_doa_mux_b0/B2_5 ;
  wire  \inst_doa_mux_b0/B2_6 ;
  wire  \inst_doa_mux_b0/B2_7 ;
  wire  \inst_doa_mux_b0/B3_0 ;
  wire  \inst_doa_mux_b0/B3_1 ;
  wire  \inst_doa_mux_b0/B3_2 ;
  wire  \inst_doa_mux_b0/B3_3 ;
  wire  \inst_doa_mux_b0/B4_0 ;
  wire  \inst_doa_mux_b0/B4_1 ;
  wire  \inst_doa_mux_b1/B0_0 ;
  wire  \inst_doa_mux_b1/B0_1 ;
  wire  \inst_doa_mux_b1/B0_10 ;
  wire  \inst_doa_mux_b1/B0_11 ;
  wire  \inst_doa_mux_b1/B0_12 ;
  wire  \inst_doa_mux_b1/B0_13 ;
  wire  \inst_doa_mux_b1/B0_14 ;
  wire  \inst_doa_mux_b1/B0_15 ;
  wire  \inst_doa_mux_b1/B0_16 ;
  wire  \inst_doa_mux_b1/B0_17 ;
  wire  \inst_doa_mux_b1/B0_18 ;
  wire  \inst_doa_mux_b1/B0_19 ;
  wire  \inst_doa_mux_b1/B0_2 ;
  wire  \inst_doa_mux_b1/B0_20 ;
  wire  \inst_doa_mux_b1/B0_21 ;
  wire  \inst_doa_mux_b1/B0_22 ;
  wire  \inst_doa_mux_b1/B0_23 ;
  wire  \inst_doa_mux_b1/B0_24 ;
  wire  \inst_doa_mux_b1/B0_25 ;
  wire  \inst_doa_mux_b1/B0_26 ;
  wire  \inst_doa_mux_b1/B0_27 ;
  wire  \inst_doa_mux_b1/B0_28 ;
  wire  \inst_doa_mux_b1/B0_29 ;
  wire  \inst_doa_mux_b1/B0_3 ;
  wire  \inst_doa_mux_b1/B0_30 ;
  wire  \inst_doa_mux_b1/B0_31 ;
  wire  \inst_doa_mux_b1/B0_4 ;
  wire  \inst_doa_mux_b1/B0_5 ;
  wire  \inst_doa_mux_b1/B0_6 ;
  wire  \inst_doa_mux_b1/B0_7 ;
  wire  \inst_doa_mux_b1/B0_8 ;
  wire  \inst_doa_mux_b1/B0_9 ;
  wire  \inst_doa_mux_b1/B1_0 ;
  wire  \inst_doa_mux_b1/B1_1 ;
  wire  \inst_doa_mux_b1/B1_10 ;
  wire  \inst_doa_mux_b1/B1_11 ;
  wire  \inst_doa_mux_b1/B1_12 ;
  wire  \inst_doa_mux_b1/B1_13 ;
  wire  \inst_doa_mux_b1/B1_14 ;
  wire  \inst_doa_mux_b1/B1_15 ;
  wire  \inst_doa_mux_b1/B1_2 ;
  wire  \inst_doa_mux_b1/B1_3 ;
  wire  \inst_doa_mux_b1/B1_4 ;
  wire  \inst_doa_mux_b1/B1_5 ;
  wire  \inst_doa_mux_b1/B1_6 ;
  wire  \inst_doa_mux_b1/B1_7 ;
  wire  \inst_doa_mux_b1/B1_8 ;
  wire  \inst_doa_mux_b1/B1_9 ;
  wire  \inst_doa_mux_b1/B2_0 ;
  wire  \inst_doa_mux_b1/B2_1 ;
  wire  \inst_doa_mux_b1/B2_2 ;
  wire  \inst_doa_mux_b1/B2_3 ;
  wire  \inst_doa_mux_b1/B2_4 ;
  wire  \inst_doa_mux_b1/B2_5 ;
  wire  \inst_doa_mux_b1/B2_6 ;
  wire  \inst_doa_mux_b1/B2_7 ;
  wire  \inst_doa_mux_b1/B3_0 ;
  wire  \inst_doa_mux_b1/B3_1 ;
  wire  \inst_doa_mux_b1/B3_2 ;
  wire  \inst_doa_mux_b1/B3_3 ;
  wire  \inst_doa_mux_b1/B4_0 ;
  wire  \inst_doa_mux_b1/B4_1 ;
  wire  \inst_doa_mux_b10/B3_0 ;
  wire  \inst_doa_mux_b10/B3_1 ;
  wire  \inst_doa_mux_b10/B3_2 ;
  wire  \inst_doa_mux_b10/B3_3 ;
  wire  \inst_doa_mux_b10/B4_0 ;
  wire  \inst_doa_mux_b10/B4_1 ;
  wire  \inst_doa_mux_b11/B3_0 ;
  wire  \inst_doa_mux_b11/B3_1 ;
  wire  \inst_doa_mux_b11/B3_2 ;
  wire  \inst_doa_mux_b11/B3_3 ;
  wire  \inst_doa_mux_b11/B4_0 ;
  wire  \inst_doa_mux_b11/B4_1 ;
  wire  \inst_doa_mux_b2/B0_0 ;
  wire  \inst_doa_mux_b2/B0_1 ;
  wire  \inst_doa_mux_b2/B0_10 ;
  wire  \inst_doa_mux_b2/B0_11 ;
  wire  \inst_doa_mux_b2/B0_12 ;
  wire  \inst_doa_mux_b2/B0_13 ;
  wire  \inst_doa_mux_b2/B0_14 ;
  wire  \inst_doa_mux_b2/B0_15 ;
  wire  \inst_doa_mux_b2/B0_16 ;
  wire  \inst_doa_mux_b2/B0_17 ;
  wire  \inst_doa_mux_b2/B0_18 ;
  wire  \inst_doa_mux_b2/B0_19 ;
  wire  \inst_doa_mux_b2/B0_2 ;
  wire  \inst_doa_mux_b2/B0_20 ;
  wire  \inst_doa_mux_b2/B0_21 ;
  wire  \inst_doa_mux_b2/B0_22 ;
  wire  \inst_doa_mux_b2/B0_23 ;
  wire  \inst_doa_mux_b2/B0_24 ;
  wire  \inst_doa_mux_b2/B0_25 ;
  wire  \inst_doa_mux_b2/B0_26 ;
  wire  \inst_doa_mux_b2/B0_27 ;
  wire  \inst_doa_mux_b2/B0_28 ;
  wire  \inst_doa_mux_b2/B0_29 ;
  wire  \inst_doa_mux_b2/B0_3 ;
  wire  \inst_doa_mux_b2/B0_30 ;
  wire  \inst_doa_mux_b2/B0_31 ;
  wire  \inst_doa_mux_b2/B0_4 ;
  wire  \inst_doa_mux_b2/B0_5 ;
  wire  \inst_doa_mux_b2/B0_6 ;
  wire  \inst_doa_mux_b2/B0_7 ;
  wire  \inst_doa_mux_b2/B0_8 ;
  wire  \inst_doa_mux_b2/B0_9 ;
  wire  \inst_doa_mux_b2/B1_0 ;
  wire  \inst_doa_mux_b2/B1_1 ;
  wire  \inst_doa_mux_b2/B1_10 ;
  wire  \inst_doa_mux_b2/B1_11 ;
  wire  \inst_doa_mux_b2/B1_12 ;
  wire  \inst_doa_mux_b2/B1_13 ;
  wire  \inst_doa_mux_b2/B1_14 ;
  wire  \inst_doa_mux_b2/B1_15 ;
  wire  \inst_doa_mux_b2/B1_2 ;
  wire  \inst_doa_mux_b2/B1_3 ;
  wire  \inst_doa_mux_b2/B1_4 ;
  wire  \inst_doa_mux_b2/B1_5 ;
  wire  \inst_doa_mux_b2/B1_6 ;
  wire  \inst_doa_mux_b2/B1_7 ;
  wire  \inst_doa_mux_b2/B1_8 ;
  wire  \inst_doa_mux_b2/B1_9 ;
  wire  \inst_doa_mux_b2/B2_0 ;
  wire  \inst_doa_mux_b2/B2_1 ;
  wire  \inst_doa_mux_b2/B2_2 ;
  wire  \inst_doa_mux_b2/B2_3 ;
  wire  \inst_doa_mux_b2/B2_4 ;
  wire  \inst_doa_mux_b2/B2_5 ;
  wire  \inst_doa_mux_b2/B2_6 ;
  wire  \inst_doa_mux_b2/B2_7 ;
  wire  \inst_doa_mux_b2/B3_0 ;
  wire  \inst_doa_mux_b2/B3_1 ;
  wire  \inst_doa_mux_b2/B3_2 ;
  wire  \inst_doa_mux_b2/B3_3 ;
  wire  \inst_doa_mux_b2/B4_0 ;
  wire  \inst_doa_mux_b2/B4_1 ;
  wire  \inst_doa_mux_b3/B0_0 ;
  wire  \inst_doa_mux_b3/B0_1 ;
  wire  \inst_doa_mux_b3/B0_10 ;
  wire  \inst_doa_mux_b3/B0_11 ;
  wire  \inst_doa_mux_b3/B0_12 ;
  wire  \inst_doa_mux_b3/B0_13 ;
  wire  \inst_doa_mux_b3/B0_14 ;
  wire  \inst_doa_mux_b3/B0_15 ;
  wire  \inst_doa_mux_b3/B0_16 ;
  wire  \inst_doa_mux_b3/B0_17 ;
  wire  \inst_doa_mux_b3/B0_18 ;
  wire  \inst_doa_mux_b3/B0_19 ;
  wire  \inst_doa_mux_b3/B0_2 ;
  wire  \inst_doa_mux_b3/B0_20 ;
  wire  \inst_doa_mux_b3/B0_21 ;
  wire  \inst_doa_mux_b3/B0_22 ;
  wire  \inst_doa_mux_b3/B0_23 ;
  wire  \inst_doa_mux_b3/B0_24 ;
  wire  \inst_doa_mux_b3/B0_25 ;
  wire  \inst_doa_mux_b3/B0_26 ;
  wire  \inst_doa_mux_b3/B0_27 ;
  wire  \inst_doa_mux_b3/B0_28 ;
  wire  \inst_doa_mux_b3/B0_29 ;
  wire  \inst_doa_mux_b3/B0_3 ;
  wire  \inst_doa_mux_b3/B0_30 ;
  wire  \inst_doa_mux_b3/B0_31 ;
  wire  \inst_doa_mux_b3/B0_4 ;
  wire  \inst_doa_mux_b3/B0_5 ;
  wire  \inst_doa_mux_b3/B0_6 ;
  wire  \inst_doa_mux_b3/B0_7 ;
  wire  \inst_doa_mux_b3/B0_8 ;
  wire  \inst_doa_mux_b3/B0_9 ;
  wire  \inst_doa_mux_b3/B1_0 ;
  wire  \inst_doa_mux_b3/B1_1 ;
  wire  \inst_doa_mux_b3/B1_10 ;
  wire  \inst_doa_mux_b3/B1_11 ;
  wire  \inst_doa_mux_b3/B1_12 ;
  wire  \inst_doa_mux_b3/B1_13 ;
  wire  \inst_doa_mux_b3/B1_14 ;
  wire  \inst_doa_mux_b3/B1_15 ;
  wire  \inst_doa_mux_b3/B1_2 ;
  wire  \inst_doa_mux_b3/B1_3 ;
  wire  \inst_doa_mux_b3/B1_4 ;
  wire  \inst_doa_mux_b3/B1_5 ;
  wire  \inst_doa_mux_b3/B1_6 ;
  wire  \inst_doa_mux_b3/B1_7 ;
  wire  \inst_doa_mux_b3/B1_8 ;
  wire  \inst_doa_mux_b3/B1_9 ;
  wire  \inst_doa_mux_b3/B2_0 ;
  wire  \inst_doa_mux_b3/B2_1 ;
  wire  \inst_doa_mux_b3/B2_2 ;
  wire  \inst_doa_mux_b3/B2_3 ;
  wire  \inst_doa_mux_b3/B2_4 ;
  wire  \inst_doa_mux_b3/B2_5 ;
  wire  \inst_doa_mux_b3/B2_6 ;
  wire  \inst_doa_mux_b3/B2_7 ;
  wire  \inst_doa_mux_b3/B3_0 ;
  wire  \inst_doa_mux_b3/B3_1 ;
  wire  \inst_doa_mux_b3/B3_2 ;
  wire  \inst_doa_mux_b3/B3_3 ;
  wire  \inst_doa_mux_b3/B4_0 ;
  wire  \inst_doa_mux_b3/B4_1 ;
  wire  \inst_doa_mux_b4/B0_0 ;
  wire  \inst_doa_mux_b4/B0_1 ;
  wire  \inst_doa_mux_b4/B0_10 ;
  wire  \inst_doa_mux_b4/B0_11 ;
  wire  \inst_doa_mux_b4/B0_12 ;
  wire  \inst_doa_mux_b4/B0_13 ;
  wire  \inst_doa_mux_b4/B0_14 ;
  wire  \inst_doa_mux_b4/B0_15 ;
  wire  \inst_doa_mux_b4/B0_16 ;
  wire  \inst_doa_mux_b4/B0_17 ;
  wire  \inst_doa_mux_b4/B0_18 ;
  wire  \inst_doa_mux_b4/B0_19 ;
  wire  \inst_doa_mux_b4/B0_2 ;
  wire  \inst_doa_mux_b4/B0_20 ;
  wire  \inst_doa_mux_b4/B0_21 ;
  wire  \inst_doa_mux_b4/B0_22 ;
  wire  \inst_doa_mux_b4/B0_23 ;
  wire  \inst_doa_mux_b4/B0_24 ;
  wire  \inst_doa_mux_b4/B0_25 ;
  wire  \inst_doa_mux_b4/B0_26 ;
  wire  \inst_doa_mux_b4/B0_27 ;
  wire  \inst_doa_mux_b4/B0_28 ;
  wire  \inst_doa_mux_b4/B0_29 ;
  wire  \inst_doa_mux_b4/B0_3 ;
  wire  \inst_doa_mux_b4/B0_30 ;
  wire  \inst_doa_mux_b4/B0_31 ;
  wire  \inst_doa_mux_b4/B0_4 ;
  wire  \inst_doa_mux_b4/B0_5 ;
  wire  \inst_doa_mux_b4/B0_6 ;
  wire  \inst_doa_mux_b4/B0_7 ;
  wire  \inst_doa_mux_b4/B0_8 ;
  wire  \inst_doa_mux_b4/B0_9 ;
  wire  \inst_doa_mux_b4/B1_0 ;
  wire  \inst_doa_mux_b4/B1_1 ;
  wire  \inst_doa_mux_b4/B1_10 ;
  wire  \inst_doa_mux_b4/B1_11 ;
  wire  \inst_doa_mux_b4/B1_12 ;
  wire  \inst_doa_mux_b4/B1_13 ;
  wire  \inst_doa_mux_b4/B1_14 ;
  wire  \inst_doa_mux_b4/B1_15 ;
  wire  \inst_doa_mux_b4/B1_2 ;
  wire  \inst_doa_mux_b4/B1_3 ;
  wire  \inst_doa_mux_b4/B1_4 ;
  wire  \inst_doa_mux_b4/B1_5 ;
  wire  \inst_doa_mux_b4/B1_6 ;
  wire  \inst_doa_mux_b4/B1_7 ;
  wire  \inst_doa_mux_b4/B1_8 ;
  wire  \inst_doa_mux_b4/B1_9 ;
  wire  \inst_doa_mux_b4/B2_0 ;
  wire  \inst_doa_mux_b4/B2_1 ;
  wire  \inst_doa_mux_b4/B2_2 ;
  wire  \inst_doa_mux_b4/B2_3 ;
  wire  \inst_doa_mux_b4/B2_4 ;
  wire  \inst_doa_mux_b4/B2_5 ;
  wire  \inst_doa_mux_b4/B2_6 ;
  wire  \inst_doa_mux_b4/B2_7 ;
  wire  \inst_doa_mux_b4/B3_0 ;
  wire  \inst_doa_mux_b4/B3_1 ;
  wire  \inst_doa_mux_b4/B3_2 ;
  wire  \inst_doa_mux_b4/B3_3 ;
  wire  \inst_doa_mux_b4/B4_0 ;
  wire  \inst_doa_mux_b4/B4_1 ;
  wire  \inst_doa_mux_b5/B0_0 ;
  wire  \inst_doa_mux_b5/B0_1 ;
  wire  \inst_doa_mux_b5/B0_10 ;
  wire  \inst_doa_mux_b5/B0_11 ;
  wire  \inst_doa_mux_b5/B0_12 ;
  wire  \inst_doa_mux_b5/B0_13 ;
  wire  \inst_doa_mux_b5/B0_14 ;
  wire  \inst_doa_mux_b5/B0_15 ;
  wire  \inst_doa_mux_b5/B0_16 ;
  wire  \inst_doa_mux_b5/B0_17 ;
  wire  \inst_doa_mux_b5/B0_18 ;
  wire  \inst_doa_mux_b5/B0_19 ;
  wire  \inst_doa_mux_b5/B0_2 ;
  wire  \inst_doa_mux_b5/B0_20 ;
  wire  \inst_doa_mux_b5/B0_21 ;
  wire  \inst_doa_mux_b5/B0_22 ;
  wire  \inst_doa_mux_b5/B0_23 ;
  wire  \inst_doa_mux_b5/B0_24 ;
  wire  \inst_doa_mux_b5/B0_25 ;
  wire  \inst_doa_mux_b5/B0_26 ;
  wire  \inst_doa_mux_b5/B0_27 ;
  wire  \inst_doa_mux_b5/B0_28 ;
  wire  \inst_doa_mux_b5/B0_29 ;
  wire  \inst_doa_mux_b5/B0_3 ;
  wire  \inst_doa_mux_b5/B0_30 ;
  wire  \inst_doa_mux_b5/B0_31 ;
  wire  \inst_doa_mux_b5/B0_4 ;
  wire  \inst_doa_mux_b5/B0_5 ;
  wire  \inst_doa_mux_b5/B0_6 ;
  wire  \inst_doa_mux_b5/B0_7 ;
  wire  \inst_doa_mux_b5/B0_8 ;
  wire  \inst_doa_mux_b5/B0_9 ;
  wire  \inst_doa_mux_b5/B1_0 ;
  wire  \inst_doa_mux_b5/B1_1 ;
  wire  \inst_doa_mux_b5/B1_10 ;
  wire  \inst_doa_mux_b5/B1_11 ;
  wire  \inst_doa_mux_b5/B1_12 ;
  wire  \inst_doa_mux_b5/B1_13 ;
  wire  \inst_doa_mux_b5/B1_14 ;
  wire  \inst_doa_mux_b5/B1_15 ;
  wire  \inst_doa_mux_b5/B1_2 ;
  wire  \inst_doa_mux_b5/B1_3 ;
  wire  \inst_doa_mux_b5/B1_4 ;
  wire  \inst_doa_mux_b5/B1_5 ;
  wire  \inst_doa_mux_b5/B1_6 ;
  wire  \inst_doa_mux_b5/B1_7 ;
  wire  \inst_doa_mux_b5/B1_8 ;
  wire  \inst_doa_mux_b5/B1_9 ;
  wire  \inst_doa_mux_b5/B2_0 ;
  wire  \inst_doa_mux_b5/B2_1 ;
  wire  \inst_doa_mux_b5/B2_2 ;
  wire  \inst_doa_mux_b5/B2_3 ;
  wire  \inst_doa_mux_b5/B2_4 ;
  wire  \inst_doa_mux_b5/B2_5 ;
  wire  \inst_doa_mux_b5/B2_6 ;
  wire  \inst_doa_mux_b5/B2_7 ;
  wire  \inst_doa_mux_b5/B3_0 ;
  wire  \inst_doa_mux_b5/B3_1 ;
  wire  \inst_doa_mux_b5/B3_2 ;
  wire  \inst_doa_mux_b5/B3_3 ;
  wire  \inst_doa_mux_b5/B4_0 ;
  wire  \inst_doa_mux_b5/B4_1 ;
  wire  \inst_doa_mux_b6/B0_0 ;
  wire  \inst_doa_mux_b6/B0_1 ;
  wire  \inst_doa_mux_b6/B0_10 ;
  wire  \inst_doa_mux_b6/B0_11 ;
  wire  \inst_doa_mux_b6/B0_12 ;
  wire  \inst_doa_mux_b6/B0_13 ;
  wire  \inst_doa_mux_b6/B0_14 ;
  wire  \inst_doa_mux_b6/B0_15 ;
  wire  \inst_doa_mux_b6/B0_16 ;
  wire  \inst_doa_mux_b6/B0_17 ;
  wire  \inst_doa_mux_b6/B0_18 ;
  wire  \inst_doa_mux_b6/B0_19 ;
  wire  \inst_doa_mux_b6/B0_2 ;
  wire  \inst_doa_mux_b6/B0_20 ;
  wire  \inst_doa_mux_b6/B0_21 ;
  wire  \inst_doa_mux_b6/B0_22 ;
  wire  \inst_doa_mux_b6/B0_23 ;
  wire  \inst_doa_mux_b6/B0_24 ;
  wire  \inst_doa_mux_b6/B0_25 ;
  wire  \inst_doa_mux_b6/B0_26 ;
  wire  \inst_doa_mux_b6/B0_27 ;
  wire  \inst_doa_mux_b6/B0_28 ;
  wire  \inst_doa_mux_b6/B0_29 ;
  wire  \inst_doa_mux_b6/B0_3 ;
  wire  \inst_doa_mux_b6/B0_30 ;
  wire  \inst_doa_mux_b6/B0_31 ;
  wire  \inst_doa_mux_b6/B0_4 ;
  wire  \inst_doa_mux_b6/B0_5 ;
  wire  \inst_doa_mux_b6/B0_6 ;
  wire  \inst_doa_mux_b6/B0_7 ;
  wire  \inst_doa_mux_b6/B0_8 ;
  wire  \inst_doa_mux_b6/B0_9 ;
  wire  \inst_doa_mux_b6/B1_0 ;
  wire  \inst_doa_mux_b6/B1_1 ;
  wire  \inst_doa_mux_b6/B1_10 ;
  wire  \inst_doa_mux_b6/B1_11 ;
  wire  \inst_doa_mux_b6/B1_12 ;
  wire  \inst_doa_mux_b6/B1_13 ;
  wire  \inst_doa_mux_b6/B1_14 ;
  wire  \inst_doa_mux_b6/B1_15 ;
  wire  \inst_doa_mux_b6/B1_2 ;
  wire  \inst_doa_mux_b6/B1_3 ;
  wire  \inst_doa_mux_b6/B1_4 ;
  wire  \inst_doa_mux_b6/B1_5 ;
  wire  \inst_doa_mux_b6/B1_6 ;
  wire  \inst_doa_mux_b6/B1_7 ;
  wire  \inst_doa_mux_b6/B1_8 ;
  wire  \inst_doa_mux_b6/B1_9 ;
  wire  \inst_doa_mux_b6/B2_0 ;
  wire  \inst_doa_mux_b6/B2_1 ;
  wire  \inst_doa_mux_b6/B2_2 ;
  wire  \inst_doa_mux_b6/B2_3 ;
  wire  \inst_doa_mux_b6/B2_4 ;
  wire  \inst_doa_mux_b6/B2_5 ;
  wire  \inst_doa_mux_b6/B2_6 ;
  wire  \inst_doa_mux_b6/B2_7 ;
  wire  \inst_doa_mux_b6/B3_0 ;
  wire  \inst_doa_mux_b6/B3_1 ;
  wire  \inst_doa_mux_b6/B3_2 ;
  wire  \inst_doa_mux_b6/B3_3 ;
  wire  \inst_doa_mux_b6/B4_0 ;
  wire  \inst_doa_mux_b6/B4_1 ;
  wire  \inst_doa_mux_b7/B0_0 ;
  wire  \inst_doa_mux_b7/B0_1 ;
  wire  \inst_doa_mux_b7/B0_10 ;
  wire  \inst_doa_mux_b7/B0_11 ;
  wire  \inst_doa_mux_b7/B0_12 ;
  wire  \inst_doa_mux_b7/B0_13 ;
  wire  \inst_doa_mux_b7/B0_14 ;
  wire  \inst_doa_mux_b7/B0_15 ;
  wire  \inst_doa_mux_b7/B0_16 ;
  wire  \inst_doa_mux_b7/B0_17 ;
  wire  \inst_doa_mux_b7/B0_18 ;
  wire  \inst_doa_mux_b7/B0_19 ;
  wire  \inst_doa_mux_b7/B0_2 ;
  wire  \inst_doa_mux_b7/B0_20 ;
  wire  \inst_doa_mux_b7/B0_21 ;
  wire  \inst_doa_mux_b7/B0_22 ;
  wire  \inst_doa_mux_b7/B0_23 ;
  wire  \inst_doa_mux_b7/B0_24 ;
  wire  \inst_doa_mux_b7/B0_25 ;
  wire  \inst_doa_mux_b7/B0_26 ;
  wire  \inst_doa_mux_b7/B0_27 ;
  wire  \inst_doa_mux_b7/B0_28 ;
  wire  \inst_doa_mux_b7/B0_29 ;
  wire  \inst_doa_mux_b7/B0_3 ;
  wire  \inst_doa_mux_b7/B0_30 ;
  wire  \inst_doa_mux_b7/B0_31 ;
  wire  \inst_doa_mux_b7/B0_4 ;
  wire  \inst_doa_mux_b7/B0_5 ;
  wire  \inst_doa_mux_b7/B0_6 ;
  wire  \inst_doa_mux_b7/B0_7 ;
  wire  \inst_doa_mux_b7/B0_8 ;
  wire  \inst_doa_mux_b7/B0_9 ;
  wire  \inst_doa_mux_b7/B1_0 ;
  wire  \inst_doa_mux_b7/B1_1 ;
  wire  \inst_doa_mux_b7/B1_10 ;
  wire  \inst_doa_mux_b7/B1_11 ;
  wire  \inst_doa_mux_b7/B1_12 ;
  wire  \inst_doa_mux_b7/B1_13 ;
  wire  \inst_doa_mux_b7/B1_14 ;
  wire  \inst_doa_mux_b7/B1_15 ;
  wire  \inst_doa_mux_b7/B1_2 ;
  wire  \inst_doa_mux_b7/B1_3 ;
  wire  \inst_doa_mux_b7/B1_4 ;
  wire  \inst_doa_mux_b7/B1_5 ;
  wire  \inst_doa_mux_b7/B1_6 ;
  wire  \inst_doa_mux_b7/B1_7 ;
  wire  \inst_doa_mux_b7/B1_8 ;
  wire  \inst_doa_mux_b7/B1_9 ;
  wire  \inst_doa_mux_b7/B2_0 ;
  wire  \inst_doa_mux_b7/B2_1 ;
  wire  \inst_doa_mux_b7/B2_2 ;
  wire  \inst_doa_mux_b7/B2_3 ;
  wire  \inst_doa_mux_b7/B2_4 ;
  wire  \inst_doa_mux_b7/B2_5 ;
  wire  \inst_doa_mux_b7/B2_6 ;
  wire  \inst_doa_mux_b7/B2_7 ;
  wire  \inst_doa_mux_b7/B3_0 ;
  wire  \inst_doa_mux_b7/B3_1 ;
  wire  \inst_doa_mux_b7/B3_2 ;
  wire  \inst_doa_mux_b7/B3_3 ;
  wire  \inst_doa_mux_b7/B4_0 ;
  wire  \inst_doa_mux_b7/B4_1 ;
  wire  \inst_doa_mux_b8/B0_0 ;
  wire  \inst_doa_mux_b8/B0_1 ;
  wire  \inst_doa_mux_b8/B0_10 ;
  wire  \inst_doa_mux_b8/B0_11 ;
  wire  \inst_doa_mux_b8/B0_12 ;
  wire  \inst_doa_mux_b8/B0_13 ;
  wire  \inst_doa_mux_b8/B0_14 ;
  wire  \inst_doa_mux_b8/B0_15 ;
  wire  \inst_doa_mux_b8/B0_16 ;
  wire  \inst_doa_mux_b8/B0_17 ;
  wire  \inst_doa_mux_b8/B0_18 ;
  wire  \inst_doa_mux_b8/B0_19 ;
  wire  \inst_doa_mux_b8/B0_2 ;
  wire  \inst_doa_mux_b8/B0_20 ;
  wire  \inst_doa_mux_b8/B0_21 ;
  wire  \inst_doa_mux_b8/B0_22 ;
  wire  \inst_doa_mux_b8/B0_23 ;
  wire  \inst_doa_mux_b8/B0_24 ;
  wire  \inst_doa_mux_b8/B0_25 ;
  wire  \inst_doa_mux_b8/B0_26 ;
  wire  \inst_doa_mux_b8/B0_27 ;
  wire  \inst_doa_mux_b8/B0_28 ;
  wire  \inst_doa_mux_b8/B0_29 ;
  wire  \inst_doa_mux_b8/B0_3 ;
  wire  \inst_doa_mux_b8/B0_30 ;
  wire  \inst_doa_mux_b8/B0_31 ;
  wire  \inst_doa_mux_b8/B0_4 ;
  wire  \inst_doa_mux_b8/B0_5 ;
  wire  \inst_doa_mux_b8/B0_6 ;
  wire  \inst_doa_mux_b8/B0_7 ;
  wire  \inst_doa_mux_b8/B0_8 ;
  wire  \inst_doa_mux_b8/B0_9 ;
  wire  \inst_doa_mux_b8/B1_0 ;
  wire  \inst_doa_mux_b8/B1_1 ;
  wire  \inst_doa_mux_b8/B1_10 ;
  wire  \inst_doa_mux_b8/B1_11 ;
  wire  \inst_doa_mux_b8/B1_12 ;
  wire  \inst_doa_mux_b8/B1_13 ;
  wire  \inst_doa_mux_b8/B1_14 ;
  wire  \inst_doa_mux_b8/B1_15 ;
  wire  \inst_doa_mux_b8/B1_2 ;
  wire  \inst_doa_mux_b8/B1_3 ;
  wire  \inst_doa_mux_b8/B1_4 ;
  wire  \inst_doa_mux_b8/B1_5 ;
  wire  \inst_doa_mux_b8/B1_6 ;
  wire  \inst_doa_mux_b8/B1_7 ;
  wire  \inst_doa_mux_b8/B1_8 ;
  wire  \inst_doa_mux_b8/B1_9 ;
  wire  \inst_doa_mux_b8/B2_0 ;
  wire  \inst_doa_mux_b8/B2_1 ;
  wire  \inst_doa_mux_b8/B2_2 ;
  wire  \inst_doa_mux_b8/B2_3 ;
  wire  \inst_doa_mux_b8/B2_4 ;
  wire  \inst_doa_mux_b8/B2_5 ;
  wire  \inst_doa_mux_b8/B2_6 ;
  wire  \inst_doa_mux_b8/B2_7 ;
  wire  \inst_doa_mux_b8/B3_0 ;
  wire  \inst_doa_mux_b8/B3_1 ;
  wire  \inst_doa_mux_b8/B3_2 ;
  wire  \inst_doa_mux_b8/B3_3 ;
  wire  \inst_doa_mux_b8/B4_0 ;
  wire  \inst_doa_mux_b8/B4_1 ;
  wire  \inst_doa_mux_b9/B3_0 ;
  wire  \inst_doa_mux_b9/B3_1 ;
  wire  \inst_doa_mux_b9/B3_2 ;
  wire  \inst_doa_mux_b9/B3_3 ;
  wire  \inst_doa_mux_b9/B4_0 ;
  wire  \inst_doa_mux_b9/B4_1 ;
  wire \and_Naddra[12]_Naddr_o ;
  wire \and_Naddra[12]_Naddr_o_al_n28 ;
  wire \and_Naddra[12]_Naddr_o_al_n60 ;
  wire \and_Naddra[12]_Naddr_o_al_n92 ;
  wire \and_Naddra[12]_addra_o ;
  wire \and_Naddra[12]_addra_o_al_n108 ;
  wire \and_Naddra[12]_addra_o_al_n44 ;
  wire \and_Naddra[12]_addra_o_al_n76 ;
  wire \and_addra[12]_Naddra_o ;
  wire \and_addra[12]_Naddra_o_al_n100 ;
  wire \and_addra[12]_Naddra_o_al_n36 ;
  wire \and_addra[12]_Naddra_o_al_n68 ;
  wire \and_addra[12]_addra[_o ;
  wire \and_addra[12]_addra[_o_al_n116 ;
  wire \and_addra[12]_addra[_o_al_n52 ;
  wire \and_addra[12]_addra[_o_al_n84 ;
  wire inst_doa_i0_000;
  wire inst_doa_i0_001;
  wire inst_doa_i0_002;
  wire inst_doa_i0_003;
  wire inst_doa_i0_004;
  wire inst_doa_i0_005;
  wire inst_doa_i0_006;
  wire inst_doa_i0_007;
  wire inst_doa_i0_008;
  wire inst_doa_i0_009;
  wire inst_doa_i0_010;
  wire inst_doa_i10_000;
  wire inst_doa_i10_001;
  wire inst_doa_i10_002;
  wire inst_doa_i10_003;
  wire inst_doa_i10_004;
  wire inst_doa_i10_005;
  wire inst_doa_i10_006;
  wire inst_doa_i10_007;
  wire inst_doa_i10_008;
  wire inst_doa_i11_000;
  wire inst_doa_i11_001;
  wire inst_doa_i11_002;
  wire inst_doa_i11_003;
  wire inst_doa_i11_004;
  wire inst_doa_i11_005;
  wire inst_doa_i11_006;
  wire inst_doa_i11_007;
  wire inst_doa_i11_008;
  wire inst_doa_i12_000;
  wire inst_doa_i12_001;
  wire inst_doa_i12_002;
  wire inst_doa_i12_003;
  wire inst_doa_i12_004;
  wire inst_doa_i12_005;
  wire inst_doa_i12_006;
  wire inst_doa_i12_007;
  wire inst_doa_i12_008;
  wire inst_doa_i13_000;
  wire inst_doa_i13_001;
  wire inst_doa_i13_002;
  wire inst_doa_i13_003;
  wire inst_doa_i13_004;
  wire inst_doa_i13_005;
  wire inst_doa_i13_006;
  wire inst_doa_i13_007;
  wire inst_doa_i13_008;
  wire inst_doa_i14_000;
  wire inst_doa_i14_001;
  wire inst_doa_i14_002;
  wire inst_doa_i14_003;
  wire inst_doa_i14_004;
  wire inst_doa_i14_005;
  wire inst_doa_i14_006;
  wire inst_doa_i14_007;
  wire inst_doa_i14_008;
  wire inst_doa_i15_000;
  wire inst_doa_i15_001;
  wire inst_doa_i15_002;
  wire inst_doa_i15_003;
  wire inst_doa_i15_004;
  wire inst_doa_i15_005;
  wire inst_doa_i15_006;
  wire inst_doa_i15_007;
  wire inst_doa_i15_008;
  wire inst_doa_i16_000;
  wire inst_doa_i16_001;
  wire inst_doa_i16_002;
  wire inst_doa_i16_003;
  wire inst_doa_i16_004;
  wire inst_doa_i16_005;
  wire inst_doa_i16_006;
  wire inst_doa_i16_007;
  wire inst_doa_i16_008;
  wire inst_doa_i16_009;
  wire inst_doa_i16_010;
  wire inst_doa_i16_011;
  wire inst_doa_i17_000;
  wire inst_doa_i17_001;
  wire inst_doa_i17_002;
  wire inst_doa_i17_003;
  wire inst_doa_i17_004;
  wire inst_doa_i17_005;
  wire inst_doa_i17_006;
  wire inst_doa_i17_007;
  wire inst_doa_i17_008;
  wire inst_doa_i18_000;
  wire inst_doa_i18_001;
  wire inst_doa_i18_002;
  wire inst_doa_i18_003;
  wire inst_doa_i18_004;
  wire inst_doa_i18_005;
  wire inst_doa_i18_006;
  wire inst_doa_i18_007;
  wire inst_doa_i18_008;
  wire inst_doa_i19_000;
  wire inst_doa_i19_001;
  wire inst_doa_i19_002;
  wire inst_doa_i19_003;
  wire inst_doa_i19_004;
  wire inst_doa_i19_005;
  wire inst_doa_i19_006;
  wire inst_doa_i19_007;
  wire inst_doa_i19_008;
  wire inst_doa_i1_000;
  wire inst_doa_i1_001;
  wire inst_doa_i1_002;
  wire inst_doa_i1_003;
  wire inst_doa_i1_004;
  wire inst_doa_i1_005;
  wire inst_doa_i1_006;
  wire inst_doa_i1_007;
  wire inst_doa_i1_008;
  wire inst_doa_i20_000;
  wire inst_doa_i20_001;
  wire inst_doa_i20_002;
  wire inst_doa_i20_003;
  wire inst_doa_i20_004;
  wire inst_doa_i20_005;
  wire inst_doa_i20_006;
  wire inst_doa_i20_007;
  wire inst_doa_i20_008;
  wire inst_doa_i21_000;
  wire inst_doa_i21_001;
  wire inst_doa_i21_002;
  wire inst_doa_i21_003;
  wire inst_doa_i21_004;
  wire inst_doa_i21_005;
  wire inst_doa_i21_006;
  wire inst_doa_i21_007;
  wire inst_doa_i21_008;
  wire inst_doa_i22_000;
  wire inst_doa_i22_001;
  wire inst_doa_i22_002;
  wire inst_doa_i22_003;
  wire inst_doa_i22_004;
  wire inst_doa_i22_005;
  wire inst_doa_i22_006;
  wire inst_doa_i22_007;
  wire inst_doa_i22_008;
  wire inst_doa_i23_000;
  wire inst_doa_i23_001;
  wire inst_doa_i23_002;
  wire inst_doa_i23_003;
  wire inst_doa_i23_004;
  wire inst_doa_i23_005;
  wire inst_doa_i23_006;
  wire inst_doa_i23_007;
  wire inst_doa_i23_008;
  wire inst_doa_i24_000;
  wire inst_doa_i24_001;
  wire inst_doa_i24_002;
  wire inst_doa_i24_003;
  wire inst_doa_i24_004;
  wire inst_doa_i24_005;
  wire inst_doa_i24_006;
  wire inst_doa_i24_007;
  wire inst_doa_i24_008;
  wire inst_doa_i24_009;
  wire inst_doa_i24_010;
  wire inst_doa_i25_000;
  wire inst_doa_i25_001;
  wire inst_doa_i25_002;
  wire inst_doa_i25_003;
  wire inst_doa_i25_004;
  wire inst_doa_i25_005;
  wire inst_doa_i25_006;
  wire inst_doa_i25_007;
  wire inst_doa_i25_008;
  wire inst_doa_i26_000;
  wire inst_doa_i26_001;
  wire inst_doa_i26_002;
  wire inst_doa_i26_003;
  wire inst_doa_i26_004;
  wire inst_doa_i26_005;
  wire inst_doa_i26_006;
  wire inst_doa_i26_007;
  wire inst_doa_i26_008;
  wire inst_doa_i27_000;
  wire inst_doa_i27_001;
  wire inst_doa_i27_002;
  wire inst_doa_i27_003;
  wire inst_doa_i27_004;
  wire inst_doa_i27_005;
  wire inst_doa_i27_006;
  wire inst_doa_i27_007;
  wire inst_doa_i27_008;
  wire inst_doa_i28_000;
  wire inst_doa_i28_001;
  wire inst_doa_i28_002;
  wire inst_doa_i28_003;
  wire inst_doa_i28_004;
  wire inst_doa_i28_005;
  wire inst_doa_i28_006;
  wire inst_doa_i28_007;
  wire inst_doa_i28_008;
  wire inst_doa_i29_000;
  wire inst_doa_i29_001;
  wire inst_doa_i29_002;
  wire inst_doa_i29_003;
  wire inst_doa_i29_004;
  wire inst_doa_i29_005;
  wire inst_doa_i29_006;
  wire inst_doa_i29_007;
  wire inst_doa_i29_008;
  wire inst_doa_i2_000;
  wire inst_doa_i2_001;
  wire inst_doa_i2_002;
  wire inst_doa_i2_003;
  wire inst_doa_i2_004;
  wire inst_doa_i2_005;
  wire inst_doa_i2_006;
  wire inst_doa_i2_007;
  wire inst_doa_i2_008;
  wire inst_doa_i30_000;
  wire inst_doa_i30_001;
  wire inst_doa_i30_002;
  wire inst_doa_i30_003;
  wire inst_doa_i30_004;
  wire inst_doa_i30_005;
  wire inst_doa_i30_006;
  wire inst_doa_i30_007;
  wire inst_doa_i30_008;
  wire inst_doa_i31_000;
  wire inst_doa_i31_001;
  wire inst_doa_i31_002;
  wire inst_doa_i31_003;
  wire inst_doa_i31_004;
  wire inst_doa_i31_005;
  wire inst_doa_i31_006;
  wire inst_doa_i31_007;
  wire inst_doa_i31_008;
  wire inst_doa_i32_000;
  wire inst_doa_i32_001;
  wire inst_doa_i32_002;
  wire inst_doa_i32_003;
  wire inst_doa_i32_004;
  wire inst_doa_i32_005;
  wire inst_doa_i32_006;
  wire inst_doa_i32_007;
  wire inst_doa_i32_008;
  wire inst_doa_i32_009;
  wire inst_doa_i32_010;
  wire inst_doa_i33_000;
  wire inst_doa_i33_001;
  wire inst_doa_i33_002;
  wire inst_doa_i33_003;
  wire inst_doa_i33_004;
  wire inst_doa_i33_005;
  wire inst_doa_i33_006;
  wire inst_doa_i33_007;
  wire inst_doa_i33_008;
  wire inst_doa_i34_000;
  wire inst_doa_i34_001;
  wire inst_doa_i34_002;
  wire inst_doa_i34_003;
  wire inst_doa_i34_004;
  wire inst_doa_i34_005;
  wire inst_doa_i34_006;
  wire inst_doa_i34_007;
  wire inst_doa_i34_008;
  wire inst_doa_i35_000;
  wire inst_doa_i35_001;
  wire inst_doa_i35_002;
  wire inst_doa_i35_003;
  wire inst_doa_i35_004;
  wire inst_doa_i35_005;
  wire inst_doa_i35_006;
  wire inst_doa_i35_007;
  wire inst_doa_i35_008;
  wire inst_doa_i36_000;
  wire inst_doa_i36_001;
  wire inst_doa_i36_002;
  wire inst_doa_i36_003;
  wire inst_doa_i36_004;
  wire inst_doa_i36_005;
  wire inst_doa_i36_006;
  wire inst_doa_i36_007;
  wire inst_doa_i36_008;
  wire inst_doa_i37_000;
  wire inst_doa_i37_001;
  wire inst_doa_i37_002;
  wire inst_doa_i37_003;
  wire inst_doa_i37_004;
  wire inst_doa_i37_005;
  wire inst_doa_i37_006;
  wire inst_doa_i37_007;
  wire inst_doa_i37_008;
  wire inst_doa_i38_000;
  wire inst_doa_i38_001;
  wire inst_doa_i38_002;
  wire inst_doa_i38_003;
  wire inst_doa_i38_004;
  wire inst_doa_i38_005;
  wire inst_doa_i38_006;
  wire inst_doa_i38_007;
  wire inst_doa_i38_008;
  wire inst_doa_i39_000;
  wire inst_doa_i39_001;
  wire inst_doa_i39_002;
  wire inst_doa_i39_003;
  wire inst_doa_i39_004;
  wire inst_doa_i39_005;
  wire inst_doa_i39_006;
  wire inst_doa_i39_007;
  wire inst_doa_i39_008;
  wire inst_doa_i3_000;
  wire inst_doa_i3_001;
  wire inst_doa_i3_002;
  wire inst_doa_i3_003;
  wire inst_doa_i3_004;
  wire inst_doa_i3_005;
  wire inst_doa_i3_006;
  wire inst_doa_i3_007;
  wire inst_doa_i3_008;
  wire inst_doa_i40_000;
  wire inst_doa_i40_001;
  wire inst_doa_i40_002;
  wire inst_doa_i40_003;
  wire inst_doa_i40_004;
  wire inst_doa_i40_005;
  wire inst_doa_i40_006;
  wire inst_doa_i40_007;
  wire inst_doa_i40_008;
  wire inst_doa_i40_009;
  wire inst_doa_i40_010;
  wire inst_doa_i40_011;
  wire inst_doa_i41_000;
  wire inst_doa_i41_001;
  wire inst_doa_i41_002;
  wire inst_doa_i41_003;
  wire inst_doa_i41_004;
  wire inst_doa_i41_005;
  wire inst_doa_i41_006;
  wire inst_doa_i41_007;
  wire inst_doa_i41_008;
  wire inst_doa_i42_000;
  wire inst_doa_i42_001;
  wire inst_doa_i42_002;
  wire inst_doa_i42_003;
  wire inst_doa_i42_004;
  wire inst_doa_i42_005;
  wire inst_doa_i42_006;
  wire inst_doa_i42_007;
  wire inst_doa_i42_008;
  wire inst_doa_i43_000;
  wire inst_doa_i43_001;
  wire inst_doa_i43_002;
  wire inst_doa_i43_003;
  wire inst_doa_i43_004;
  wire inst_doa_i43_005;
  wire inst_doa_i43_006;
  wire inst_doa_i43_007;
  wire inst_doa_i43_008;
  wire inst_doa_i44_000;
  wire inst_doa_i44_001;
  wire inst_doa_i44_002;
  wire inst_doa_i44_003;
  wire inst_doa_i44_004;
  wire inst_doa_i44_005;
  wire inst_doa_i44_006;
  wire inst_doa_i44_007;
  wire inst_doa_i44_008;
  wire inst_doa_i45_000;
  wire inst_doa_i45_001;
  wire inst_doa_i45_002;
  wire inst_doa_i45_003;
  wire inst_doa_i45_004;
  wire inst_doa_i45_005;
  wire inst_doa_i45_006;
  wire inst_doa_i45_007;
  wire inst_doa_i45_008;
  wire inst_doa_i46_000;
  wire inst_doa_i46_001;
  wire inst_doa_i46_002;
  wire inst_doa_i46_003;
  wire inst_doa_i46_004;
  wire inst_doa_i46_005;
  wire inst_doa_i46_006;
  wire inst_doa_i46_007;
  wire inst_doa_i46_008;
  wire inst_doa_i47_000;
  wire inst_doa_i47_001;
  wire inst_doa_i47_002;
  wire inst_doa_i47_003;
  wire inst_doa_i47_004;
  wire inst_doa_i47_005;
  wire inst_doa_i47_006;
  wire inst_doa_i47_007;
  wire inst_doa_i47_008;
  wire inst_doa_i48_000;
  wire inst_doa_i48_001;
  wire inst_doa_i48_002;
  wire inst_doa_i48_003;
  wire inst_doa_i48_004;
  wire inst_doa_i48_005;
  wire inst_doa_i48_006;
  wire inst_doa_i48_007;
  wire inst_doa_i48_008;
  wire inst_doa_i48_009;
  wire inst_doa_i48_010;
  wire inst_doa_i48_011;
  wire inst_doa_i49_000;
  wire inst_doa_i49_001;
  wire inst_doa_i49_002;
  wire inst_doa_i49_003;
  wire inst_doa_i49_004;
  wire inst_doa_i49_005;
  wire inst_doa_i49_006;
  wire inst_doa_i49_007;
  wire inst_doa_i49_008;
  wire inst_doa_i4_000;
  wire inst_doa_i4_001;
  wire inst_doa_i4_002;
  wire inst_doa_i4_003;
  wire inst_doa_i4_004;
  wire inst_doa_i4_005;
  wire inst_doa_i4_006;
  wire inst_doa_i4_007;
  wire inst_doa_i4_008;
  wire inst_doa_i50_000;
  wire inst_doa_i50_001;
  wire inst_doa_i50_002;
  wire inst_doa_i50_003;
  wire inst_doa_i50_004;
  wire inst_doa_i50_005;
  wire inst_doa_i50_006;
  wire inst_doa_i50_007;
  wire inst_doa_i50_008;
  wire inst_doa_i51_000;
  wire inst_doa_i51_001;
  wire inst_doa_i51_002;
  wire inst_doa_i51_003;
  wire inst_doa_i51_004;
  wire inst_doa_i51_005;
  wire inst_doa_i51_006;
  wire inst_doa_i51_007;
  wire inst_doa_i51_008;
  wire inst_doa_i52_000;
  wire inst_doa_i52_001;
  wire inst_doa_i52_002;
  wire inst_doa_i52_003;
  wire inst_doa_i52_004;
  wire inst_doa_i52_005;
  wire inst_doa_i52_006;
  wire inst_doa_i52_007;
  wire inst_doa_i52_008;
  wire inst_doa_i53_000;
  wire inst_doa_i53_001;
  wire inst_doa_i53_002;
  wire inst_doa_i53_003;
  wire inst_doa_i53_004;
  wire inst_doa_i53_005;
  wire inst_doa_i53_006;
  wire inst_doa_i53_007;
  wire inst_doa_i53_008;
  wire inst_doa_i54_000;
  wire inst_doa_i54_001;
  wire inst_doa_i54_002;
  wire inst_doa_i54_003;
  wire inst_doa_i54_004;
  wire inst_doa_i54_005;
  wire inst_doa_i54_006;
  wire inst_doa_i54_007;
  wire inst_doa_i54_008;
  wire inst_doa_i55_000;
  wire inst_doa_i55_001;
  wire inst_doa_i55_002;
  wire inst_doa_i55_003;
  wire inst_doa_i55_004;
  wire inst_doa_i55_005;
  wire inst_doa_i55_006;
  wire inst_doa_i55_007;
  wire inst_doa_i55_008;
  wire inst_doa_i56_000;
  wire inst_doa_i56_001;
  wire inst_doa_i56_002;
  wire inst_doa_i56_003;
  wire inst_doa_i56_004;
  wire inst_doa_i56_005;
  wire inst_doa_i56_006;
  wire inst_doa_i56_007;
  wire inst_doa_i56_008;
  wire inst_doa_i56_009;
  wire inst_doa_i56_010;
  wire inst_doa_i57_000;
  wire inst_doa_i57_001;
  wire inst_doa_i57_002;
  wire inst_doa_i57_003;
  wire inst_doa_i57_004;
  wire inst_doa_i57_005;
  wire inst_doa_i57_006;
  wire inst_doa_i57_007;
  wire inst_doa_i57_008;
  wire inst_doa_i58_000;
  wire inst_doa_i58_001;
  wire inst_doa_i58_002;
  wire inst_doa_i58_003;
  wire inst_doa_i58_004;
  wire inst_doa_i58_005;
  wire inst_doa_i58_006;
  wire inst_doa_i58_007;
  wire inst_doa_i58_008;
  wire inst_doa_i59_000;
  wire inst_doa_i59_001;
  wire inst_doa_i59_002;
  wire inst_doa_i59_003;
  wire inst_doa_i59_004;
  wire inst_doa_i59_005;
  wire inst_doa_i59_006;
  wire inst_doa_i59_007;
  wire inst_doa_i59_008;
  wire inst_doa_i5_000;
  wire inst_doa_i5_001;
  wire inst_doa_i5_002;
  wire inst_doa_i5_003;
  wire inst_doa_i5_004;
  wire inst_doa_i5_005;
  wire inst_doa_i5_006;
  wire inst_doa_i5_007;
  wire inst_doa_i5_008;
  wire inst_doa_i60_000;
  wire inst_doa_i60_001;
  wire inst_doa_i60_002;
  wire inst_doa_i60_003;
  wire inst_doa_i60_004;
  wire inst_doa_i60_005;
  wire inst_doa_i60_006;
  wire inst_doa_i60_007;
  wire inst_doa_i60_008;
  wire inst_doa_i61_000;
  wire inst_doa_i61_001;
  wire inst_doa_i61_002;
  wire inst_doa_i61_003;
  wire inst_doa_i61_004;
  wire inst_doa_i61_005;
  wire inst_doa_i61_006;
  wire inst_doa_i61_007;
  wire inst_doa_i61_008;
  wire inst_doa_i62_000;
  wire inst_doa_i62_001;
  wire inst_doa_i62_002;
  wire inst_doa_i62_003;
  wire inst_doa_i62_004;
  wire inst_doa_i62_005;
  wire inst_doa_i62_006;
  wire inst_doa_i62_007;
  wire inst_doa_i62_008;
  wire inst_doa_i63_000;
  wire inst_doa_i63_001;
  wire inst_doa_i63_002;
  wire inst_doa_i63_003;
  wire inst_doa_i63_004;
  wire inst_doa_i63_005;
  wire inst_doa_i63_006;
  wire inst_doa_i63_007;
  wire inst_doa_i63_008;
  wire inst_doa_i6_000;
  wire inst_doa_i6_001;
  wire inst_doa_i6_002;
  wire inst_doa_i6_003;
  wire inst_doa_i6_004;
  wire inst_doa_i6_005;
  wire inst_doa_i6_006;
  wire inst_doa_i6_007;
  wire inst_doa_i6_008;
  wire inst_doa_i7_000;
  wire inst_doa_i7_001;
  wire inst_doa_i7_002;
  wire inst_doa_i7_003;
  wire inst_doa_i7_004;
  wire inst_doa_i7_005;
  wire inst_doa_i7_006;
  wire inst_doa_i7_007;
  wire inst_doa_i7_008;
  wire inst_doa_i8_000;
  wire inst_doa_i8_001;
  wire inst_doa_i8_002;
  wire inst_doa_i8_003;
  wire inst_doa_i8_004;
  wire inst_doa_i8_005;
  wire inst_doa_i8_006;
  wire inst_doa_i8_007;
  wire inst_doa_i8_008;
  wire inst_doa_i8_009;
  wire inst_doa_i8_010;
  wire inst_doa_i8_011;
  wire inst_doa_i9_000;
  wire inst_doa_i9_001;
  wire inst_doa_i9_002;
  wire inst_doa_i9_003;
  wire inst_doa_i9_004;
  wire inst_doa_i9_005;
  wire inst_doa_i9_006;
  wire inst_doa_i9_007;
  wire inst_doa_i9_008;

  AL_DFF_X addra_pipe_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clka),
    .d(addra[10]),
    .en(1'b1),
    .sr(rsta),
    .ss(1'b0),
    .q(addra_piped[0]));
  AL_DFF_X addra_pipe_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clka),
    .d(addra[11]),
    .en(1'b1),
    .sr(rsta),
    .ss(1'b0),
    .q(addra_piped[1]));
  AL_DFF_X addra_pipe_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clka),
    .d(addra[12]),
    .en(1'b1),
    .sr(rsta),
    .ss(1'b0),
    .q(addra_piped[2]));
  AL_DFF_X addra_pipe_b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clka),
    .d(addra[13]),
    .en(1'b1),
    .sr(rsta),
    .ss(1'b0),
    .q(addra_piped[3]));
  AL_DFF_X addra_pipe_b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clka),
    .d(addra[14]),
    .en(1'b1),
    .sr(rsta),
    .ss(1'b0),
    .q(addra_piped[4]));
  AL_DFF_X addra_pipe_b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clka),
    .d(addra[15]),
    .en(1'b1),
    .sr(rsta),
    .ss(1'b0),
    .q(addra_piped[5]));
  and \and_Naddra[12]_Naddr  (\and_Naddra[12]_Naddr_o , ~addra[12], ~addra[13], ~addra[14], ~addra[15]);
  and \and_Naddra[12]_Naddr_al_u28  (\and_Naddra[12]_Naddr_o_al_n28 , ~addra[12], ~addra[13], addra[14], ~addra[15]);
  and \and_Naddra[12]_Naddr_al_u60  (\and_Naddra[12]_Naddr_o_al_n60 , ~addra[12], ~addra[13], ~addra[14], addra[15]);
  and \and_Naddra[12]_Naddr_al_u92  (\and_Naddra[12]_Naddr_o_al_n92 , ~addra[12], ~addra[13], addra[14], addra[15]);
  and \and_Naddra[12]_addra  (\and_Naddra[12]_addra_o , ~addra[12], addra[13], ~addra[14], ~addra[15]);
  and \and_Naddra[12]_addra_al_u108  (\and_Naddra[12]_addra_o_al_n108 , ~addra[12], addra[13], addra[14], addra[15]);
  and \and_Naddra[12]_addra_al_u44  (\and_Naddra[12]_addra_o_al_n44 , ~addra[12], addra[13], addra[14], ~addra[15]);
  and \and_Naddra[12]_addra_al_u76  (\and_Naddra[12]_addra_o_al_n76 , ~addra[12], addra[13], ~addra[14], addra[15]);
  and \and_addra[12]_Naddra  (\and_addra[12]_Naddra_o , addra[12], ~addra[13], ~addra[14], ~addra[15]);
  and \and_addra[12]_Naddra_al_u100  (\and_addra[12]_Naddra_o_al_n100 , addra[12], ~addra[13], addra[14], addra[15]);
  and \and_addra[12]_Naddra_al_u36  (\and_addra[12]_Naddra_o_al_n36 , addra[12], ~addra[13], addra[14], ~addra[15]);
  and \and_addra[12]_Naddra_al_u68  (\and_addra[12]_Naddra_o_al_n68 , addra[12], ~addra[13], ~addra[14], addra[15]);
  and \and_addra[12]_addra[  (\and_addra[12]_addra[_o , addra[12], addra[13], ~addra[14], ~addra[15]);
  and \and_addra[12]_addra[_al_u116  (\and_addra[12]_addra[_o_al_n116 , addra[12], addra[13], addra[14], addra[15]);
  and \and_addra[12]_addra[_al_u52  (\and_addra[12]_addra[_o_al_n52 , addra[12], addra[13], addra[14], ~addra[15]);
  and \and_addra[12]_addra[_al_u84  (\and_addra[12]_addra[_o_al_n84 , addra[12], addra[13], ~addra[14], addra[15]);
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  // address_offset=0;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFFFFFFFFFFFFFF),
    .INIT_08(256'hFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE),
    .INIT_09(256'hFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE),
    .INIT_0A(256'hFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE),
    .INIT_0B(256'hFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE),
    .INIT_0C(256'hFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE),
    .INIT_0D(256'hFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFD),
    .INIT_0E(256'hFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFD),
    .INIT_0F(256'hFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFD),
    .INIT_10(256'hFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFDFDFDFD),
    .INIT_11(256'hFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFC),
    .INIT_12(256'hFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFC),
    .INIT_13(256'hFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFCFC),
    .INIT_14(256'hFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFB),
    .INIT_15(256'hFAFAFAFAFAFAFAFAFAFAFAFAFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFB),
    .INIT_16(256'hFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFA),
    .INIT_17(256'hF9F9F9FAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFA),
    .INIT_18(256'hF9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9),
    .INIT_19(256'hF9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9),
    .INIT_1A(256'hF8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8),
    .INIT_1B(256'hF7F7F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8),
    .INIT_1C(256'hF7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7),
    .INIT_1D(256'hF6F6F6F6F6F6F6F6F6F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7),
    .INIT_1E(256'hF6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6),
    .INIT_1F(256'hF5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F6F6F6F6F6F6F6F6F6F6F6F6F6F6),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_000000_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_Naddr_o ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i0_008,inst_doa_i0_007,inst_doa_i0_006,inst_doa_i0_005,inst_doa_i0_004,inst_doa_i0_003,inst_doa_i0_002,inst_doa_i0_001,inst_doa_i0_000}));
  // address_offset=0;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'h000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_000000_009 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n108,open_n109,open_n110,open_n111,open_n112,open_n113,open_n114,1'b0,open_n115}),
    .rsta(rsta),
    .doa({open_n130,open_n131,open_n132,open_n133,open_n134,open_n135,open_n136,open_n137,inst_doa_i0_009}));
  // address_offset=0;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_000000_010 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n166,open_n167,open_n168,open_n169,open_n170,open_n171,open_n172,1'b0,open_n173}),
    .rsta(rsta),
    .doa({open_n188,open_n189,open_n190,open_n191,open_n192,open_n193,open_n194,open_n195,inst_doa_i0_010}));
  // address_offset=1024;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'hF5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5),
    .INIT_01(256'hF4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F5),
    .INIT_02(256'hF3F3F3F3F3F3F3F3F3F3F3F3F3F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4),
    .INIT_03(256'hF3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3),
    .INIT_04(256'hF2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F3F3),
    .INIT_05(256'hF1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2),
    .INIT_06(256'hF0F0F0F0F0F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1),
    .INIT_07(256'hF0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0),
    .INIT_08(256'hEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFF0F0F0F0F0),
    .INIT_09(256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEFEFEFEFEFEFEFEFEFEFEFEFEFEF),
    .INIT_0A(256'hEDEDEDEDEDEDEDEDEDEDEDEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE),
    .INIT_0B(256'hECECECECEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDED),
    .INIT_0C(256'hECECECECECECECECECECECECECECECECECECECECECECECECECECECECECECECEC),
    .INIT_0D(256'hEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEC),
    .INIT_0E(256'hEAEAEAEAEAEAEAEAEAEAEAEAEAEAEAEAEAEAEAEAEAEAEAEAEAEAEBEBEBEBEBEB),
    .INIT_0F(256'hE9E9E9E9E9E9E9E9E9E9E9E9E9E9E9E9E9E9E9E9E9E9E9EAEAEAEAEAEAEAEAEA),
    .INIT_10(256'hE8E8E8E8E8E8E8E8E8E8E8E8E8E8E8E8E8E8E8E8E9E9E9E9E9E9E9E9E9E9E9E9),
    .INIT_11(256'hE7E7E7E7E7E7E7E7E7E7E7E7E7E7E7E7E7E7E8E8E8E8E8E8E8E8E8E8E8E8E8E8),
    .INIT_12(256'hE6E6E6E6E6E6E6E6E6E6E6E6E6E6E6E6E7E7E7E7E7E7E7E7E7E7E7E7E7E7E7E7),
    .INIT_13(256'hE5E5E5E5E5E5E5E5E5E5E5E5E5E5E5E5E6E6E6E6E6E6E6E6E6E6E6E6E6E6E6E6),
    .INIT_14(256'hE4E4E4E4E4E4E4E4E4E4E4E4E4E4E4E4E5E5E5E5E5E5E5E5E5E5E5E5E5E5E5E5),
    .INIT_15(256'hE3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E4E4E4E4E4E4E4E4E4E4E4E4E4E4E4E4),
    .INIT_16(256'hE2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3),
    .INIT_17(256'hE1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E2E2E2E2E2E2E2E2E2E2E2E2E2),
    .INIT_18(256'hE0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E1E1E1E1E1E1E1E1E1E1E1),
    .INIT_19(256'hDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFE0E0E0E0E0E0E0E0),
    .INIT_1A(256'hDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDFDFDFDFDF),
    .INIT_1B(256'hDCDCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDEDE),
    .INIT_1C(256'hDBDBDBDBDBDBDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDC),
    .INIT_1D(256'hDADADADADADADADADADADADBDBDBDBDBDBDBDBDBDBDBDBDBDBDBDBDBDBDBDBDB),
    .INIT_1E(256'hD9D9D9D9D9D9D9D9D9D9D9D9D9D9D9D9DADADADADADADADADADADADADADADADA),
    .INIT_1F(256'hD8D8D8D8D8D8D8D8D8D8D8D8D8D8D8D8D8D8D8D8D8D8D9D9D9D9D9D9D9D9D9D9),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_001024_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_Naddr_o ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i1_008,inst_doa_i1_007,inst_doa_i1_006,inst_doa_i1_005,inst_doa_i1_004,inst_doa_i1_003,inst_doa_i1_002,inst_doa_i1_001,inst_doa_i1_000}));
  // address_offset=2048;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'hD6D7D7D7D7D7D7D7D7D7D7D7D7D7D7D7D7D7D7D7D7D7D7D7D7D7D7D8D8D8D8D8),
    .INIT_01(256'hD5D5D5D5D5D5D5D5D6D6D6D6D6D6D6D6D6D6D6D6D6D6D6D6D6D6D6D6D6D6D6D6),
    .INIT_02(256'hD4D4D4D4D4D4D4D4D4D4D4D4D4D4D4D5D5D5D5D5D5D5D5D5D5D5D5D5D5D5D5D5),
    .INIT_03(256'hD3D3D3D3D3D3D3D3D3D3D3D3D3D3D3D3D3D3D3D3D3D3D4D4D4D4D4D4D4D4D4D4),
    .INIT_04(256'hD1D1D1D1D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D3D3D3),
    .INIT_05(256'hD0D0D0D0D0D0D0D0D0D0D0D0D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1),
    .INIT_06(256'hCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFD0D0D0D0D0D0D0D0D0D0D0D0),
    .INIT_07(256'hCDCDCDCDCDCECECECECECECECECECECECECECECECECECECECECECECECECFCFCF),
    .INIT_08(256'hCCCCCCCCCCCCCCCCCCCCCCCCCCCCCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCD),
    .INIT_09(256'hCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCCCCCCCCCCCCCCCCCC),
    .INIT_0A(256'hC9C9C9C9C9C9C9C9C9C9CACACACACACACACACACACACACACACACACACACACACACA),
    .INIT_0B(256'hC8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C9C9C9C9C9C9C9C9C9C9C9C9),
    .INIT_0C(256'hC6C6C6C6C6C6C6C7C7C7C7C7C7C7C7C7C7C7C7C7C7C7C7C7C7C7C7C7C7C8C8C8),
    .INIT_0D(256'hC5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C6C6C6C6C6C6C6C6C6C6C6C6C6C6),
    .INIT_0E(256'hC3C3C3C3C3C3C3C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C5C5C5C5),
    .INIT_0F(256'hC2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C3C3C3C3C3C3C3C3C3C3C3C3C3C3),
    .INIT_10(256'hC0C0C0C0C0C0C0C0C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C2C2C2),
    .INIT_11(256'hBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFC0C0C0C0C0C0C0C0C0C0C0C0C0),
    .INIT_12(256'hBDBDBDBDBDBDBDBDBDBDBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBFBF),
    .INIT_13(256'hBBBBBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBDBDBDBDBDBDBDBDBDBD),
    .INIT_14(256'hBABABABABABABABABABABABABABABBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB),
    .INIT_15(256'hB8B8B8B8B8B8B9B9B9B9B9B9B9B9B9B9B9B9B9B9B9B9B9B9B9B9BABABABABABA),
    .INIT_16(256'hB7B7B7B7B7B7B7B7B7B7B7B7B7B7B7B7B7B7B7B8B8B8B8B8B8B8B8B8B8B8B8B8),
    .INIT_17(256'hB5B5B5B5B5B5B5B5B5B5B5B5B6B6B6B6B6B6B6B6B6B6B6B6B6B6B6B6B6B6B6B6),
    .INIT_18(256'hB3B3B3B3B3B3B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B5B5B5B5B5B5B5),
    .INIT_19(256'hB1B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B3B3B3B3B3B3B3B3B3B3B3B3B3),
    .INIT_1A(256'hB0B0B0B0B0B0B0B0B0B0B0B0B0B0B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1),
    .INIT_1B(256'hAEAEAEAEAEAEAEAEAEAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFB0B0B0B0B0),
    .INIT_1C(256'hACACACACACADADADADADADADADADADADADADADADADADADAEAEAEAEAEAEAEAEAE),
    .INIT_1D(256'hABABABABABABABABABABABABABABABABABABACACACACACACACACACACACACACAC),
    .INIT_1E(256'hA9A9A9A9A9A9A9A9A9A9A9A9A9A9A9AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA),
    .INIT_1F(256'hA7A7A7A7A7A7A7A7A7A7A7A8A8A8A8A8A8A8A8A8A8A8A8A8A8A8A8A8A8A9A9A9),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_002048_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_Naddr_o ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i2_008,inst_doa_i2_007,inst_doa_i2_006,inst_doa_i2_005,inst_doa_i2_004,inst_doa_i2_003,inst_doa_i2_002,inst_doa_i2_001,inst_doa_i2_000}));
  // address_offset=3072;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'hA5A5A5A5A5A5A5A5A6A6A6A6A6A6A6A6A6A6A6A6A6A6A6A6A6A6A7A7A7A7A7A7),
    .INIT_01(256'hA3A3A3A3A3A4A4A4A4A4A4A4A4A4A4A4A4A4A4A4A4A4A4A5A5A5A5A5A5A5A5A5),
    .INIT_02(256'hA1A1A1A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A3A3A3A3A3A3A3A3A3A3A3A3),
    .INIT_03(256'h9FA0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A1A1A1A1A1A1A1A1A1A1A1A1A1A1),
    .INIT_04(256'h9E9E9E9E9E9E9E9E9E9E9E9E9E9E9E9E9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F),
    .INIT_05(256'h9C9C9C9C9C9C9C9C9C9C9C9C9C9C9C9D9D9D9D9D9D9D9D9D9D9D9D9D9D9D9D9D),
    .INIT_06(256'h9A9A9A9A9A9A9A9A9A9A9A9A9A9A9B9B9B9B9B9B9B9B9B9B9B9B9B9B9B9B9C9C),
    .INIT_07(256'h9898989898989898989898989899999999999999999999999999999999999A9A),
    .INIT_08(256'h9696969696969696969696969697979797979797979797979797979797989898),
    .INIT_09(256'h9494949494949494949494949495959595959595959595959595959595969696),
    .INIT_0A(256'h9292929292929292929292929293939393939393939393939393939393949494),
    .INIT_0B(256'h9090909090909090909090909091919191919191919191919191919191929292),
    .INIT_0C(256'h8E8E8E8E8E8E8E8E8E8E8E8E8E8E8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F909090),
    .INIT_0D(256'h8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8D8D8D8D8D8D8D8D8D8D8D8D8D8D8D8E8E),
    .INIT_0E(256'h898A8A8A8A8A8A8A8A8A8A8A8A8A8A8A8B8B8B8B8B8B8B8B8B8B8B8B8B8B8B8C),
    .INIT_0F(256'h8787888888888888888888888888888888888989898989898989898989898989),
    .INIT_10(256'h8585858586868686868686868686868686868687878787878787878787878787),
    .INIT_11(256'h8383838383838484848484848484848484848484848585858585858585858585),
    .INIT_12(256'h8181818181818181818282828282828282828282828282838383838383838383),
    .INIT_13(256'h7F7F7F7F7F7F7F7F7F7F7F808080808080808080808080808080818181818181),
    .INIT_14(256'h7D7D7D7D7D7D7D7D7D7D7D7D7D7D7E7E7E7E7E7E7E7E7E7E7E7E7E7E7E7F7F7F),
    .INIT_15(256'h7A7A7A7B7B7B7B7B7B7B7B7B7B7B7B7B7B7C7C7C7C7C7C7C7C7C7C7C7C7C7C7D),
    .INIT_16(256'h78787878787879797979797979797979797979797A7A7A7A7A7A7A7A7A7A7A7A),
    .INIT_17(256'h7676767676767676767777777777777777777777777777777878787878787878),
    .INIT_18(256'h7474747474747474747474747475757575757575757575757575757676767676),
    .INIT_19(256'h7171717272727272727272727272727272737373737373737373737373737374),
    .INIT_1A(256'h6F6F6F6F6F6F6F70707070707070707070707070707171717171717171717171),
    .INIT_1B(256'h6D6D6D6D6D6D6D6D6D6D6D6D6E6E6E6E6E6E6E6E6E6E6E6E6E6F6F6F6F6F6F6F),
    .INIT_1C(256'h6A6A6A6B6B6B6B6B6B6B6B6B6B6B6B6B6C6C6C6C6C6C6C6C6C6C6C6C6C6C6D6D),
    .INIT_1D(256'h6868686868686869696969696969696969696969696A6A6A6A6A6A6A6A6A6A6A),
    .INIT_1E(256'h6666666666666666666666666767676767676767676767676767686868686868),
    .INIT_1F(256'h6363636364646464646464646464646464646565656565656565656565656566),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_003072_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_Naddr_o ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i3_008,inst_doa_i3_007,inst_doa_i3_006,inst_doa_i3_005,inst_doa_i3_004,inst_doa_i3_003,inst_doa_i3_002,inst_doa_i3_001,inst_doa_i3_000}));
  // address_offset=4096;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'h6161616161616161616162626262626262626262626262636363636363636363),
    .INIT_01(256'h5E5E5F5F5F5F5F5F5F5F5F5F5F5F5F6060606060606060606060606061616161),
    .INIT_02(256'h5C5C5C5C5C5C5C5C5D5D5D5D5D5D5D5D5D5D5D5D5D5E5E5E5E5E5E5E5E5E5E5E),
    .INIT_03(256'h595A5A5A5A5A5A5A5A5A5A5A5A5A5B5B5B5B5B5B5B5B5B5B5B5B5B5C5C5C5C5C),
    .INIT_04(256'h5757575757575758585858585858585858585858595959595959595959595959),
    .INIT_05(256'h5455555555555555555555555555565656565656565656565656575757575757),
    .INIT_06(256'h5252525252525253535353535353535353535353545454545454545454545454),
    .INIT_07(256'h4F50505050505050505050505050515151515151515151515151515252525252),
    .INIT_08(256'h4D4D4D4D4D4D4D4D4E4E4E4E4E4E4E4E4E4E4E4E4E4F4F4F4F4F4F4F4F4F4F4F),
    .INIT_09(256'h4A4A4A4B4B4B4B4B4B4B4B4B4B4B4B4C4C4C4C4C4C4C4C4C4C4C4C4C4D4D4D4D),
    .INIT_0A(256'h48484848484848484848494949494949494949494949494A4A4A4A4A4A4A4A4A),
    .INIT_0B(256'h4545454545464646464646464646464646464747474747474747474747474848),
    .INIT_0C(256'h4243434343434343434343434344444444444444444444444445454545454545),
    .INIT_0D(256'h4040404040404040404141414141414141414141414242424242424242424242),
    .INIT_0E(256'h3D3D3D3D3E3E3E3E3E3E3E3E3E3E3E3E3F3F3F3F3F3F3F3F3F3F3F3F40404040),
    .INIT_0F(256'h3B3B3B3B3B3B3B3B3B3B3B3B3C3C3C3C3C3C3C3C3C3C3C3C3D3D3D3D3D3D3D3D),
    .INIT_10(256'h3838383838383838383939393939393939393939393A3A3A3A3A3A3A3A3A3A3A),
    .INIT_11(256'h3535353535363636363636363636363636373737373737373737373737383838),
    .INIT_12(256'h3232333333333333333333333333343434343434343434343435353535353535),
    .INIT_13(256'h3030303030303030303030313131313131313131313132323232323232323232),
    .INIT_14(256'h2D2D2D2D2D2D2D2D2E2E2E2E2E2E2E2E2E2E2E2F2F2F2F2F2F2F2F2F2F2F2F30),
    .INIT_15(256'h2A2A2A2A2A2B2B2B2B2B2B2B2B2B2B2B2B2C2C2C2C2C2C2C2C2C2C2C2D2D2D2D),
    .INIT_16(256'h27272728282828282828282828282929292929292929292929292A2A2A2A2A2A),
    .INIT_17(256'h2425252525252525252525252626262626262626262626262727272727272727),
    .INIT_18(256'h2222222222222222222223232323232323232323232324242424242424242424),
    .INIT_19(256'h1F1F1F1F1F1F1F1F1F2020202020202020202020212121212121212121212122),
    .INIT_1A(256'h1C1C1C1C1C1C1C1D1D1D1D1D1D1D1D1D1D1D1E1E1E1E1E1E1E1E1E1E1E1F1F1F),
    .INIT_1B(256'h1919191919191A1A1A1A1A1A1A1A1A1A1A1B1B1B1B1B1B1B1B1B1B1B1C1C1C1C),
    .INIT_1C(256'h1616161616171717171717171717171718181818181818181818181919191919),
    .INIT_1D(256'h1313131314141414141414141414141515151515151515151515161616161616),
    .INIT_1E(256'h1010101111111111111111111111121212121212121212121213131313131313),
    .INIT_1F(256'h0D0D0E0E0E0E0E0E0E0E0E0E0E0F0F0F0F0F0F0F0F0F0F0F1010101010101010),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_004096_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_Naddra_o ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i4_008,inst_doa_i4_007,inst_doa_i4_006,inst_doa_i4_005,inst_doa_i4_004,inst_doa_i4_003,inst_doa_i4_002,inst_doa_i4_001,inst_doa_i4_000}));
  // address_offset=5120;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0A0A0B0B0B0B0B0B0B0B0B0B0B0C0C0C0C0C0C0C0C0C0C0C0D0D0D0D0D0D0D0D),
    .INIT_01(256'h07070808080808080808080808090909090909090909090A0A0A0A0A0A0A0A0A),
    .INIT_02(256'h0404050505050505050505050506060606060606060606070707070707070707),
    .INIT_03(256'h0101020202020202020202020203030303030303030303040404040404040404),
    .INIT_04(256'hFEFEFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000101010101010101),
    .INIT_05(256'hFBFBFBFCFCFCFCFCFCFCFCFCFCFDFDFDFDFDFDFDFDFDFDFDFEFEFEFEFEFEFEFE),
    .INIT_06(256'hF8F8F8F8F9F9F9F9F9F9F9F9F9F9FAFAFAFAFAFAFAFAFAFAFAFBFBFBFBFBFBFB),
    .INIT_07(256'hF5F5F5F5F5F6F6F6F6F6F6F6F6F6F6F7F7F7F7F7F7F7F7F7F7F8F8F8F8F8F8F8),
    .INIT_08(256'hF2F2F2F2F2F2F3F3F3F3F3F3F3F3F3F3F4F4F4F4F4F4F4F4F4F4F5F5F5F5F5F5),
    .INIT_09(256'hEFEFEFEFEFEFEFF0F0F0F0F0F0F0F0F0F0F1F1F1F1F1F1F1F1F1F1F2F2F2F2F2),
    .INIT_0A(256'hECECECECECECECECEDEDEDEDEDEDEDEDEDEDEEEEEEEEEEEEEEEEEEEEEEEFEFEF),
    .INIT_0B(256'hE9E9E9E9E9E9E9E9E9E9EAEAEAEAEAEAEAEAEAEAEBEBEBEBEBEBEBEBEBEBECEC),
    .INIT_0C(256'hE5E6E6E6E6E6E6E6E6E6E6E7E7E7E7E7E7E7E7E7E7E7E8E8E8E8E8E8E8E8E8E8),
    .INIT_0D(256'hE2E2E2E3E3E3E3E3E3E3E3E3E3E4E4E4E4E4E4E4E4E4E4E5E5E5E5E5E5E5E5E5),
    .INIT_0E(256'hDFDFDFDFDFE0E0E0E0E0E0E0E0E0E0E1E1E1E1E1E1E1E1E1E1E2E2E2E2E2E2E2),
    .INIT_0F(256'hDCDCDCDCDCDCDCDDDDDDDDDDDDDDDDDDDDDEDEDEDEDEDEDEDEDEDEDFDFDFDFDF),
    .INIT_10(256'hD9D9D9D9D9D9D9D9D9D9DADADADADADADADADADADBDBDBDBDBDBDBDBDBDBDCDC),
    .INIT_11(256'hD5D5D6D6D6D6D6D6D6D6D6D6D7D7D7D7D7D7D7D7D7D7D8D8D8D8D8D8D8D8D8D8),
    .INIT_12(256'hD2D2D2D2D2D3D3D3D3D3D3D3D3D3D3D4D4D4D4D4D4D4D4D4D4D5D5D5D5D5D5D5),
    .INIT_13(256'hCFCFCFCFCFCFCFCFD0D0D0D0D0D0D0D0D0D1D1D1D1D1D1D1D1D1D1D2D2D2D2D2),
    .INIT_14(256'hCBCCCCCCCCCCCCCCCCCCCCCDCDCDCDCDCDCDCDCDCECECECECECECECECECECFCF),
    .INIT_15(256'hC8C8C8C8C9C9C9C9C9C9C9C9C9C9CACACACACACACACACACBCBCBCBCBCBCBCBCB),
    .INIT_16(256'hC5C5C5C5C5C5C5C6C6C6C6C6C6C6C6C6C6C7C7C7C7C7C7C7C7C7C8C8C8C8C8C8),
    .INIT_17(256'hC1C2C2C2C2C2C2C2C2C2C2C3C3C3C3C3C3C3C3C3C4C4C4C4C4C4C4C4C4C4C5C5),
    .INIT_18(256'hBEBEBEBEBEBFBFBFBFBFBFBFBFBFC0C0C0C0C0C0C0C0C0C0C1C1C1C1C1C1C1C1),
    .INIT_19(256'hBBBBBBBBBBBBBBBBBCBCBCBCBCBCBCBCBCBCBDBDBDBDBDBDBDBDBDBEBEBEBEBE),
    .INIT_1A(256'hB7B7B8B8B8B8B8B8B8B8B8B8B9B9B9B9B9B9B9B9B9BABABABABABABABABABABB),
    .INIT_1B(256'hB4B4B4B4B4B4B5B5B5B5B5B5B5B5B5B5B6B6B6B6B6B6B6B6B6B7B7B7B7B7B7B7),
    .INIT_1C(256'hB0B1B1B1B1B1B1B1B1B1B2B2B2B2B2B2B2B2B2B2B3B3B3B3B3B3B3B3B3B4B4B4),
    .INIT_1D(256'hADADADADADAEAEAEAEAEAEAEAEAEAFAFAFAFAFAFAFAFAFAFB0B0B0B0B0B0B0B0),
    .INIT_1E(256'hAAAAAAAAAAAAAAAAAAABABABABABABABABABABACACACACACACACACACADADADAD),
    .INIT_1F(256'hA6A6A6A6A6A7A7A7A7A7A7A7A7A7A8A8A8A8A8A8A8A8A8A9A9A9A9A9A9A9A9A9),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_005120_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_Naddra_o ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i5_008,inst_doa_i5_007,inst_doa_i5_006,inst_doa_i5_005,inst_doa_i5_004,inst_doa_i5_003,inst_doa_i5_002,inst_doa_i5_001,inst_doa_i5_000}));
  // address_offset=6144;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hA3A3A3A3A3A3A3A3A3A4A4A4A4A4A4A4A4A4A5A5A5A5A5A5A5A5A5A5A6A6A6A6),
    .INIT_01(256'h9F9F9F9F9FA0A0A0A0A0A0A0A0A0A1A1A1A1A1A1A1A1A1A2A2A2A2A2A2A2A2A2),
    .INIT_02(256'h9C9C9C9C9C9C9C9C9C9C9D9D9D9D9D9D9D9D9D9E9E9E9E9E9E9E9E9E9F9F9F9F),
    .INIT_03(256'h98989898989999999999999999999A9A9A9A9A9A9A9A9A9B9B9B9B9B9B9B9B9B),
    .INIT_04(256'h9495959595959595959596969696969696969697979797979797979798989898),
    .INIT_05(256'h9191919191919192929292929292929293939393939393939494949494949494),
    .INIT_06(256'h8D8D8D8E8E8E8E8E8E8E8E8E8F8F8F8F8F8F8F8F8F9090909090909090909191),
    .INIT_07(256'h8A8A8A8A8A8A8A8A8B8B8B8B8B8B8B8B8B8C8C8C8C8C8C8C8C8C8D8D8D8D8D8D),
    .INIT_08(256'h868686868687878787878787878788888888888888888889898989898989898A),
    .INIT_09(256'h8282838383838383838383848484848484848485858585858585858586868686),
    .INIT_0A(256'h7F7F7F7F7F7F7F7F808080808080808081818181818181818182828282828282),
    .INIT_0B(256'h7B7B7B7B7B7C7C7C7C7C7C7C7C7D7D7D7D7D7D7D7D7D7E7E7E7E7E7E7E7E7E7F),
    .INIT_0C(256'h777778787878787878787879797979797979797A7A7A7A7A7A7A7A7A7B7B7B7B),
    .INIT_0D(256'h7474747474747474757575757575757575767676767676767677777777777777),
    .INIT_0E(256'h7070707070717171717171717171727272727272727272737373737373737374),
    .INIT_0F(256'h6C6C6C6D6D6D6D6D6D6D6D6D6E6E6E6E6E6E6E6E6F6F6F6F6F6F6F6F6F707070),
    .INIT_10(256'h686969696969696969696A6A6A6A6A6A6A6A6B6B6B6B6B6B6B6B6B6C6C6C6C6C),
    .INIT_11(256'h6565656565656565666666666666666667676767676767676768686868686868),
    .INIT_12(256'h6161616161616262626262626262636363636363636363646464646464646465),
    .INIT_13(256'h5D5D5D5D5E5E5E5E5E5E5E5E5F5F5F5F5F5F5F5F5F6060606060606060616161),
    .INIT_14(256'h59595A5A5A5A5A5A5A5A5A5B5B5B5B5B5B5B5B5C5C5C5C5C5C5C5C5D5D5D5D5D),
    .INIT_15(256'h5556565656565656565757575757575757575858585858585858595959595959),
    .INIT_16(256'h5252525252525252535353535353535354545454545454545455555555555555),
    .INIT_17(256'h4E4E4E4E4E4E4E4F4F4F4F4F4F4F4F5050505050505050515151515151515151),
    .INIT_18(256'h4A4A4A4A4A4A4B4B4B4B4B4B4B4B4C4C4C4C4C4C4C4C4D4D4D4D4D4D4D4D4E4E),
    .INIT_19(256'h46464646464747474747474747484848484848484849494949494949494A4A4A),
    .INIT_1A(256'h4242424243434343434343434444444444444444454545454545454546464646),
    .INIT_1B(256'h3E3E3E3F3F3F3F3F3F3F3F404040404040404041414141414141414142424242),
    .INIT_1C(256'h3A3A3A3B3B3B3B3B3B3B3B3C3C3C3C3C3C3C3C3D3D3D3D3D3D3D3D3E3E3E3E3E),
    .INIT_1D(256'h36363737373737373737383838383838383839393939393939393A3A3A3A3A3A),
    .INIT_1E(256'h3232333333333333333334343434343434343535353535353535363636363636),
    .INIT_1F(256'h2E2E2F2F2F2F2F2F2F2F30303030303030303131313131313131323232323232),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_006144_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_Naddra_o ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i6_008,inst_doa_i6_007,inst_doa_i6_006,inst_doa_i6_005,inst_doa_i6_004,inst_doa_i6_003,inst_doa_i6_002,inst_doa_i6_001,inst_doa_i6_000}));
  // address_offset=7168;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'h2A2A2B2B2B2B2B2B2B2B2C2C2C2C2C2C2C2C2D2D2D2D2D2D2D2D2E2E2E2E2E2E),
    .INIT_01(256'h26262727272727272727282828282828282829292929292929292A2A2A2A2A2A),
    .INIT_02(256'h2222232323232323232324242424242424242525252525252525262626262626),
    .INIT_03(256'h1E1E1F1F1F1F1F1F1F1F20202020202020202121212121212121222222222222),
    .INIT_04(256'h1A1A1B1B1B1B1B1B1B1B1C1C1C1C1C1C1C1C1D1D1D1D1D1D1D1D1E1E1E1E1E1E),
    .INIT_05(256'h1616161717171717171717181818181818181819191919191919191A1A1A1A1A),
    .INIT_06(256'h1212121213131313131313141414141414141415151515151515151616161616),
    .INIT_07(256'h0E0E0E0E0F0F0F0F0F0F0F0F1010101010101010111111111111111112121212),
    .INIT_08(256'h0A0A0A0A0A0B0B0B0B0B0B0B0B0C0C0C0C0C0C0C0C0D0D0D0D0D0D0D0E0E0E0E),
    .INIT_09(256'h06060606060607070707070707070808080808080808090909090909090A0A0A),
    .INIT_0A(256'h0202020202020203030303030303030404040404040404050505050505050606),
    .INIT_0B(256'hFDFEFEFEFEFEFEFEFFFFFFFFFFFFFFFF00000000000000000101010101010102),
    .INIT_0C(256'hF9F9FAFAFAFAFAFAFAFAFBFBFBFBFBFBFBFCFCFCFCFCFCFCFCFDFDFDFDFDFDFD),
    .INIT_0D(256'hF5F5F5F6F6F6F6F6F6F6F6F7F7F7F7F7F7F7F7F8F8F8F8F8F8F8F9F9F9F9F9F9),
    .INIT_0E(256'hF1F1F1F1F1F2F2F2F2F2F2F2F3F3F3F3F3F3F3F3F4F4F4F4F4F4F4F4F5F5F5F5),
    .INIT_0F(256'hEDEDEDEDEDEDEEEEEEEEEEEEEEEEEFEFEFEFEFEFEFEFF0F0F0F0F0F0F0F1F1F1),
    .INIT_10(256'hE9E9E9E9E9E9E9E9EAEAEAEAEAEAEAEAEBEBEBEBEBEBEBECECECECECECECECED),
    .INIT_11(256'hE4E4E5E5E5E5E5E5E5E5E6E6E6E6E6E6E6E7E7E7E7E7E7E7E7E8E8E8E8E8E8E8),
    .INIT_12(256'hE0E0E0E0E1E1E1E1E1E1E1E1E2E2E2E2E2E2E2E3E3E3E3E3E3E3E3E4E4E4E4E4),
    .INIT_13(256'hDCDCDCDCDCDCDDDDDDDDDDDDDDDDDEDEDEDEDEDEDEDFDFDFDFDFDFDFDFE0E0E0),
    .INIT_14(256'hD7D8D8D8D8D8D8D8D9D9D9D9D9D9D9D9DADADADADADADADBDBDBDBDBDBDBDBDC),
    .INIT_15(256'hD3D3D3D4D4D4D4D4D4D4D5D5D5D5D5D5D5D5D6D6D6D6D6D6D6D7D7D7D7D7D7D7),
    .INIT_16(256'hCFCFCFCFCFD0D0D0D0D0D0D0D0D1D1D1D1D1D1D1D2D2D2D2D2D2D2D2D3D3D3D3),
    .INIT_17(256'hCBCBCBCBCBCBCBCBCCCCCCCCCCCCCCCDCDCDCDCDCDCDCECECECECECECECECFCF),
    .INIT_18(256'hC6C6C6C7C7C7C7C7C7C7C8C8C8C8C8C8C8C8C9C9C9C9C9C9C9CACACACACACACA),
    .INIT_19(256'hC2C2C2C2C2C3C3C3C3C3C3C3C3C4C4C4C4C4C4C4C5C5C5C5C5C5C5C6C6C6C6C6),
    .INIT_1A(256'hBDBEBEBEBEBEBEBEBFBFBFBFBFBFBFC0C0C0C0C0C0C0C0C1C1C1C1C1C1C1C2C2),
    .INIT_1B(256'hB9B9B9BABABABABABABABABBBBBBBBBBBBBBBCBCBCBCBCBCBCBDBDBDBDBDBDBD),
    .INIT_1C(256'hB5B5B5B5B5B5B6B6B6B6B6B6B6B6B7B7B7B7B7B7B7B8B8B8B8B8B8B8B9B9B9B9),
    .INIT_1D(256'hB0B0B1B1B1B1B1B1B1B2B2B2B2B2B2B2B3B3B3B3B3B3B3B3B4B4B4B4B4B4B4B5),
    .INIT_1E(256'hACACACACACADADADADADADADAEAEAEAEAEAEAEAFAFAFAFAFAFAFAFB0B0B0B0B0),
    .INIT_1F(256'hA7A8A8A8A8A8A8A8A9A9A9A9A9A9A9AAAAAAAAAAAAAAAAABABABABABABABACAC),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_007168_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_Naddra_o ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i7_008,inst_doa_i7_007,inst_doa_i7_006,inst_doa_i7_005,inst_doa_i7_004,inst_doa_i7_003,inst_doa_i7_002,inst_doa_i7_001,inst_doa_i7_000}));
  // address_offset=8192;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'hA3A3A3A3A4A4A4A4A4A4A4A5A5A5A5A5A5A5A5A6A6A6A6A6A6A6A7A7A7A7A7A7),
    .INIT_01(256'h9F9F9F9F9F9F9FA0A0A0A0A0A0A0A0A1A1A1A1A1A1A1A2A2A2A2A2A2A2A3A3A3),
    .INIT_02(256'h9A9A9A9A9B9B9B9B9B9B9B9C9C9C9C9C9C9C9D9D9D9D9D9D9D9E9E9E9E9E9E9E),
    .INIT_03(256'h96969696969696979797979797979898989898989899999999999999999A9A9A),
    .INIT_04(256'h9191919192929292929292939393939393939494949494949495959595959595),
    .INIT_05(256'h8D8D8D8D8D8D8D8E8E8E8E8E8E8E8F8F8F8F8F8F8F9090909090909090919191),
    .INIT_06(256'h88888888898989898989898A8A8A8A8A8A8A8B8B8B8B8B8B8B8C8C8C8C8C8C8C),
    .INIT_07(256'h8384848484848484858585858585858686868686868687878787878787888888),
    .INIT_08(256'h7F7F7F7F7F808080808080808181818181818182828282828282838383838383),
    .INIT_09(256'h7A7A7B7B7B7B7B7B7B7C7C7C7C7C7C7C7D7D7D7D7D7D7D7E7E7E7E7E7E7E7F7F),
    .INIT_0A(256'h7676767676767777777777777778787878787878797979797979797A7A7A7A7A),
    .INIT_0B(256'h7171717272727272727273737373737373747474747474747575757575757576),
    .INIT_0C(256'h6D6D6D6D6D6D6D6E6E6E6E6E6E6E6F6F6F6F6F6F6F7070707070707071717171),
    .INIT_0D(256'h68686868696969696969696A6A6A6A6A6A6A6B6B6B6B6B6B6B6C6C6C6C6C6C6C),
    .INIT_0E(256'h6363646464646464646565656565656566666666666666676767676767686868),
    .INIT_0F(256'h5F5F5F5F5F5F6060606060606061616161616161626262626262626363636363),
    .INIT_10(256'h5A5A5A5A5B5B5B5B5B5B5B5C5C5C5C5C5C5C5D5D5D5D5D5D5D5E5E5E5E5E5E5F),
    .INIT_11(256'h55555656565656565657575757575758585858585858595959595959595A5A5A),
    .INIT_12(256'h5151515151515252525252525253535353535353545454545454545555555555),
    .INIT_13(256'h4C4C4C4C4D4D4D4D4D4D4D4E4E4E4E4E4E4E4F4F4F4F4F4F4F50505050505050),
    .INIT_14(256'h474748484848484848494949494949494A4A4A4A4A4A4A4B4B4B4B4B4B4C4C4C),
    .INIT_15(256'h4343434343434344444444444444454545454545454646464646464647474747),
    .INIT_16(256'h3E3E3E3E3E3F3F3F3F3F3F3F4040404040404041414141414141424242424242),
    .INIT_17(256'h393939393A3A3A3A3A3A3B3B3B3B3B3B3B3C3C3C3C3C3C3C3D3D3D3D3D3D3D3E),
    .INIT_18(256'h3434353535353535353636363636363637373737373738383838383838393939),
    .INIT_19(256'h2F30303030303031313131313131323232323232323333333333333434343434),
    .INIT_1A(256'h2B2B2B2B2B2B2C2C2C2C2C2C2C2D2D2D2D2D2D2E2E2E2E2E2E2E2F2F2F2F2F2F),
    .INIT_1B(256'h262626262627272727272728282828282828292929292929292A2A2A2A2A2A2B),
    .INIT_1C(256'h2121212222222222222223232323232323242424242424252525252525252626),
    .INIT_1D(256'h1C1C1D1D1D1D1D1D1D1E1E1E1E1E1E1F1F1F1F1F1F1F20202020202020212121),
    .INIT_1E(256'h17181818181818181919191919191A1A1A1A1A1A1A1B1B1B1B1B1B1C1C1C1C1C),
    .INIT_1F(256'h1313131313131314141414141415151515151515161616161616171717171717),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_008192_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_addra_o ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i8_008,inst_doa_i8_007,inst_doa_i8_006,inst_doa_i8_005,inst_doa_i8_004,inst_doa_i8_003,inst_doa_i8_002,inst_doa_i8_001,inst_doa_i8_000}));
  // address_offset=8192;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'h0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_008192_009 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n560,open_n561,open_n562,open_n563,open_n564,open_n565,open_n566,1'b0,open_n567}),
    .rsta(rsta),
    .doa({open_n582,open_n583,open_n584,open_n585,open_n586,open_n587,open_n588,open_n589,inst_doa_i8_009}));
  // address_offset=8192;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'h0000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_008192_010 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n618,open_n619,open_n620,open_n621,open_n622,open_n623,open_n624,1'b0,open_n625}),
    .rsta(rsta),
    .doa({open_n640,open_n641,open_n642,open_n643,open_n644,open_n645,open_n646,open_n647,inst_doa_i8_010}));
  // address_offset=8192;data_offset=11;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_008192_011 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n676,open_n677,open_n678,open_n679,open_n680,open_n681,open_n682,1'b0,open_n683}),
    .rsta(rsta),
    .doa({open_n698,open_n699,open_n700,open_n701,open_n702,open_n703,open_n704,open_n705,inst_doa_i8_011}));
  // address_offset=9216;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h000000000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0E0E0E0E0E0E0F0F0F0F0F0F1010101010101011111111111112121212121212),
    .INIT_01(256'h09090909090A0A0A0A0A0A0B0B0B0B0B0B0B0C0C0C0C0C0C0C0D0D0D0D0D0D0E),
    .INIT_02(256'h0404040405050505050505060606060606070707070707070808080808080909),
    .INIT_03(256'hFFFFFF0000000000000001010101010102020202020202030303030303030404),
    .INIT_04(256'hFAFAFAFBFBFBFBFBFBFCFCFCFCFCFCFCFDFDFDFDFDFDFEFEFEFEFEFEFEFFFFFF),
    .INIT_05(256'hF5F5F6F6F6F6F6F6F6F7F7F7F7F7F7F8F8F8F8F8F8F8F9F9F9F9F9F9FAFAFAFA),
    .INIT_06(256'hF0F0F1F1F1F1F1F1F2F2F2F2F2F2F2F3F3F3F3F3F3F4F4F4F4F4F4F4F5F5F5F5),
    .INIT_07(256'hEBEBECECECECECECEDEDEDEDEDEDEEEEEEEEEEEEEEEFEFEFEFEFEFF0F0F0F0F0),
    .INIT_08(256'hE6E7E7E7E7E7E7E7E8E8E8E8E8E8E9E9E9E9E9E9E9EAEAEAEAEAEAEBEBEBEBEB),
    .INIT_09(256'hE1E2E2E2E2E2E2E3E3E3E3E3E3E3E4E4E4E4E4E4E5E5E5E5E5E5E5E6E6E6E6E6),
    .INIT_0A(256'hDCDDDDDDDDDDDDDEDEDEDEDEDEDEDFDFDFDFDFDFE0E0E0E0E0E0E0E1E1E1E1E1),
    .INIT_0B(256'hD7D8D8D8D8D8D8D9D9D9D9D9D9D9DADADADADADADBDBDBDBDBDBDBDCDCDCDCDC),
    .INIT_0C(256'hD2D3D3D3D3D3D3D4D4D4D4D4D4D4D5D5D5D5D5D5D6D6D6D6D6D6D7D7D7D7D7D7),
    .INIT_0D(256'hCDCECECECECECECFCFCFCFCFCFCFD0D0D0D0D0D0D1D1D1D1D1D1D1D2D2D2D2D2),
    .INIT_0E(256'hC8C9C9C9C9C9C9C9CACACACACACACBCBCBCBCBCBCCCCCCCCCCCCCCCDCDCDCDCD),
    .INIT_0F(256'hC3C4C4C4C4C4C4C4C5C5C5C5C5C5C6C6C6C6C6C6C7C7C7C7C7C7C7C8C8C8C8C8),
    .INIT_10(256'hBEBEBFBFBFBFBFBFC0C0C0C0C0C0C1C1C1C1C1C1C1C2C2C2C2C2C2C3C3C3C3C3),
    .INIT_11(256'hB9B9BABABABABABABBBBBBBBBBBBBBBCBCBCBCBCBCBDBDBDBDBDBDBEBEBEBEBE),
    .INIT_12(256'hB4B4B4B5B5B5B5B5B5B6B6B6B6B6B6B7B7B7B7B7B7B7B8B8B8B8B8B8B9B9B9B9),
    .INIT_13(256'hAFAFAFB0B0B0B0B0B0B1B1B1B1B1B1B1B2B2B2B2B2B2B3B3B3B3B3B3B4B4B4B4),
    .INIT_14(256'hAAAAAAAAABABABABABABACACACACACACADADADADADADADAEAEAEAEAEAEAFAFAF),
    .INIT_15(256'hA5A5A5A5A6A6A6A6A6A6A6A7A7A7A7A7A7A8A8A8A8A8A8A9A9A9A9A9A9AAAAAA),
    .INIT_16(256'hA0A0A0A0A0A1A1A1A1A1A1A2A2A2A2A2A2A2A3A3A3A3A3A3A4A4A4A4A4A4A5A5),
    .INIT_17(256'h9B9B9B9B9B9B9C9C9C9C9C9C9D9D9D9D9D9D9E9E9E9E9E9E9E9F9F9F9F9F9FA0),
    .INIT_18(256'h959696969696969797979797979898989898989999999999999A9A9A9A9A9A9A),
    .INIT_19(256'h9090919191919191929292929292939393939393949494949494959595959595),
    .INIT_1A(256'h8B8B8B8C8C8C8C8C8C8D8D8D8D8D8D8E8E8E8E8E8E8F8F8F8F8F8F9090909090),
    .INIT_1B(256'h868686868787878787878888888888888989898989898A8A8A8A8A8A8B8B8B8B),
    .INIT_1C(256'h8181818181828282828282838383838383848484848484858585858585868686),
    .INIT_1D(256'h7C7C7C7C7C7C7D7D7D7D7D7D7E7E7E7E7E7E7F7F7F7F7F7F8080808080808081),
    .INIT_1E(256'h767777777777777878787878787979797979797A7A7A7A7A7A7A7B7B7B7B7B7B),
    .INIT_1F(256'h7171727272727272727373737373737474747474747575757575757676767676),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_009216_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_addra_o ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i9_008,inst_doa_i9_007,inst_doa_i9_006,inst_doa_i9_005,inst_doa_i9_004,inst_doa_i9_003,inst_doa_i9_002,inst_doa_i9_001,inst_doa_i9_000}));
  // address_offset=10240;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'h6C6C6C6C6D6D6D6D6D6D6E6E6E6E6E6E6F6F6F6F6F6F70707070707071717171),
    .INIT_01(256'h67676767676868686868686969696969696A6A6A6A6A6A6A6B6B6B6B6B6B6C6C),
    .INIT_02(256'h6162626262626263636363636364646464646465656565656566666666666667),
    .INIT_03(256'h5C5C5D5D5D5D5D5D5E5E5E5E5E5E5F5F5F5F5F5F606060606060606161616161),
    .INIT_04(256'h575757575858585858585959595959595A5A5A5A5A5A5B5B5B5B5B5B5C5C5C5C),
    .INIT_05(256'h5252525252525353535353535454545454545555555555555656565656565757),
    .INIT_06(256'h4C4D4D4D4D4D4D4E4E4E4E4E4E4F4F4F4F4F4F50505050505051515151515152),
    .INIT_07(256'h4747474848484848484949494949494A4A4A4A4A4A4B4B4B4B4B4B4C4C4C4C4C),
    .INIT_08(256'h4242424242434343434343444444444444454545454545464646464646474747),
    .INIT_09(256'h3C3D3D3D3D3D3D3E3E3E3E3E3E3F3F3F3F3F3F40404040404041414141414142),
    .INIT_0A(256'h3737373838383838383939393939393A3A3A3A3A3A3B3B3B3B3B3B3C3C3C3C3C),
    .INIT_0B(256'h3232323232333333333333343434343434353535353535363636363636373737),
    .INIT_0C(256'h2C2D2D2D2D2D2D2E2E2E2E2E2E2F2F2F2F2F2F30303030303031313131313132),
    .INIT_0D(256'h2727272828282828282929292929292A2A2A2A2A2A2B2B2B2B2B2B2C2C2C2C2C),
    .INIT_0E(256'h2222222222232323232323242424242424252525252525262626262626272727),
    .INIT_0F(256'h1C1C1D1D1D1D1D1D1E1E1E1E1E1E1F1F1F1F1F1F202020202020212121212122),
    .INIT_10(256'h171717171818181818181919191919191A1A1A1A1A1A1B1B1B1B1B1B1C1C1C1C),
    .INIT_11(256'h1112121212121313131313131414141414141515151515151616161616161717),
    .INIT_12(256'h0C0C0C0D0D0D0D0D0D0E0E0E0E0E0E0F0F0F0F0F0F1010101010101111111111),
    .INIT_13(256'h07070707070808080808080909090909090A0A0A0A0A0A0B0B0B0B0B0B0C0C0C),
    .INIT_14(256'h0101020202020202030303030303040404040404050505050505060606060606),
    .INIT_15(256'hFCFCFCFCFCFDFDFDFDFDFDFEFEFEFEFEFFFFFFFFFFFF00000000000001010101),
    .INIT_16(256'hF6F7F7F7F7F7F7F8F8F8F8F8F8F9F9F9F9F9F9FAFAFAFAFAFAFBFBFBFBFBFBFC),
    .INIT_17(256'hF1F1F1F1F2F2F2F2F2F2F3F3F3F3F3F3F4F4F4F4F4F4F5F5F5F5F5F5F6F6F6F6),
    .INIT_18(256'hEBECECECECECECEDEDEDEDEDEDEEEEEEEEEEEEEFEFEFEFEFF0F0F0F0F0F0F1F1),
    .INIT_19(256'hE6E6E6E6E7E7E7E7E7E7E8E8E8E8E8E8E9E9E9E9E9EAEAEAEAEAEAEBEBEBEBEB),
    .INIT_1A(256'hE0E1E1E1E1E1E1E2E2E2E2E2E3E3E3E3E3E3E4E4E4E4E4E4E5E5E5E5E5E5E6E6),
    .INIT_1B(256'hDBDBDBDBDCDCDCDCDCDCDDDDDDDDDDDEDEDEDEDEDEDFDFDFDFDFDFE0E0E0E0E0),
    .INIT_1C(256'hD5D6D6D6D6D6D6D7D7D7D7D7D8D8D8D8D8D8D9D9D9D9D9D9DADADADADADADBDB),
    .INIT_1D(256'hD0D0D0D0D1D1D1D1D1D1D2D2D2D2D2D3D3D3D3D3D3D4D4D4D4D4D4D5D5D5D5D5),
    .INIT_1E(256'hCACBCBCBCBCBCBCCCCCCCCCCCCCDCDCDCDCDCECECECECECECFCFCFCFCFCFD0D0),
    .INIT_1F(256'hC5C5C5C5C6C6C6C6C6C6C7C7C7C7C7C7C8C8C8C8C8C8C9C9C9C9C9CACACACACA),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_010240_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_addra_o ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i10_008,inst_doa_i10_007,inst_doa_i10_006,inst_doa_i10_005,inst_doa_i10_004,inst_doa_i10_003,inst_doa_i10_002,inst_doa_i10_001,inst_doa_i10_000}));
  // address_offset=11264;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'hBFBFC0C0C0C0C0C1C1C1C1C1C1C2C2C2C2C2C2C3C3C3C3C3C3C4C4C4C4C4C5C5),
    .INIT_01(256'hBABABABABABBBBBBBBBBBBBCBCBCBCBCBDBDBDBDBDBDBEBEBEBEBEBEBFBFBFBF),
    .INIT_02(256'hB4B4B5B5B5B5B5B5B6B6B6B6B6B6B7B7B7B7B7B8B8B8B8B8B8B9B9B9B9B9B9BA),
    .INIT_03(256'hAFAFAFAFAFAFB0B0B0B0B0B1B1B1B1B1B1B2B2B2B2B2B2B3B3B3B3B3B4B4B4B4),
    .INIT_04(256'hA9A9A9AAAAAAAAAAAAABABABABABABACACACACACADADADADADADAEAEAEAEAEAE),
    .INIT_05(256'hA3A4A4A4A4A4A5A5A5A5A5A5A6A6A6A6A6A6A7A7A7A7A7A7A8A8A8A8A8A9A9A9),
    .INIT_06(256'h9E9E9E9E9F9F9F9F9F9FA0A0A0A0A0A0A1A1A1A1A1A2A2A2A2A2A2A3A3A3A3A3),
    .INIT_07(256'h98989999999999999A9A9A9A9A9B9B9B9B9B9B9C9C9C9C9C9C9D9D9D9D9D9E9E),
    .INIT_08(256'h9393939393949494949494959595959595969696969697979797979798989898),
    .INIT_09(256'h8D8D8D8E8E8E8E8E8E8F8F8F8F8F8F9090909090919191919191929292929292),
    .INIT_0A(256'h878888888888888989898989898A8A8A8A8A8B8B8B8B8B8B8C8C8C8C8C8C8D8D),
    .INIT_0B(256'h8282828282838383838384848484848485858585858586868686868787878787),
    .INIT_0C(256'h7C7C7C7D7D7D7D7D7E7E7E7E7E7E7F7F7F7F7F7F808080808081818181818182),
    .INIT_0D(256'h7677777777777778787878787979797979797A7A7A7A7A7B7B7B7B7B7B7C7C7C),
    .INIT_0E(256'h7171717171727272727273737373737374747474747475757575757676767676),
    .INIT_0F(256'h6B6B6B6C6C6C6C6C6D6D6D6D6D6D6E6E6E6E6E6E6F6F6F6F6F70707070707071),
    .INIT_10(256'h6566666666666667676767676868686868686969696969696A6A6A6A6A6B6B6B),
    .INIT_11(256'h6060606060616161616162626262626263636363636364646464646565656565),
    .INIT_12(256'h5A5A5A5B5B5B5B5B5B5C5C5C5C5C5D5D5D5D5D5D5E5E5E5E5E5E5F5F5F5F5F60),
    .INIT_13(256'h5454555555555556565656565657575757575858585858585959595959595A5A),
    .INIT_14(256'h4F4F4F4F4F4F5050505050515151515151525252525253535353535354545454),
    .INIT_15(256'h494949494A4A4A4A4A4A4B4B4B4B4B4C4C4C4C4C4C4D4D4D4D4D4E4E4E4E4E4E),
    .INIT_16(256'h4343444444444444454545454545464646464647474747474748484848484949),
    .INIT_17(256'h3D3E3E3E3E3E3E3F3F3F3F3F4040404040404141414141424242424242434343),
    .INIT_18(256'h38383838383939393939393A3A3A3A3A3B3B3B3B3B3B3C3C3C3C3C3D3D3D3D3D),
    .INIT_19(256'h3232323233333333333434343434343535353535363636363636373737373737),
    .INIT_1A(256'h2C2C2D2D2D2D2D2D2E2E2E2E2E2E2F2F2F2F2F30303030303031313131313232),
    .INIT_1B(256'h2627272727272728282828282929292929292A2A2A2A2A2B2B2B2B2B2B2C2C2C),
    .INIT_1C(256'h2121212121222222222222232323232323242424242425252525252526262626),
    .INIT_1D(256'h1B1B1B1B1C1C1C1C1C1C1D1D1D1D1D1E1E1E1E1E1E1F1F1F1F1F202020202020),
    .INIT_1E(256'h151515161616161616171717171718181818181819191919191A1A1A1A1A1A1B),
    .INIT_1F(256'h0F0F101010101010111111111112121212121213131313131414141414141515),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_011264_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_addra_o ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i11_008,inst_doa_i11_007,inst_doa_i11_006,inst_doa_i11_005,inst_doa_i11_004,inst_doa_i11_003,inst_doa_i11_002,inst_doa_i11_001,inst_doa_i11_000}));
  // address_offset=12288;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h090A0A0A0A0A0B0B0B0B0B0B0C0C0C0C0C0D0D0D0D0D0D0E0E0E0E0E0F0F0F0F),
    .INIT_01(256'h0404040404050505050505060606060607070707070708080808080909090909),
    .INIT_02(256'hFEFEFEFEFFFFFFFFFFFF00000000000101010101010202020202030303030303),
    .INIT_03(256'hF8F8F8F9F9F9F9F9F9FAFAFAFAFAFBFBFBFBFBFBFCFCFCFCFCFDFDFDFDFDFDFE),
    .INIT_04(256'hF2F2F2F3F3F3F3F3F4F4F4F4F4F4F5F5F5F5F5F6F6F6F6F6F6F7F7F7F7F7F8F8),
    .INIT_05(256'hECECEDEDEDEDEDEEEEEEEEEEEEEFEFEFEFEFF0F0F0F0F0F0F1F1F1F1F1F2F2F2),
    .INIT_06(256'hE6E7E7E7E7E7E8E8E8E8E8E8E9E9E9E9E9EAEAEAEAEAEAEBEBEBEBEBECECECEC),
    .INIT_07(256'hE1E1E1E1E1E1E2E2E2E2E2E3E3E3E3E3E3E4E4E4E4E4E5E5E5E5E5E6E6E6E6E6),
    .INIT_08(256'hDBDBDBDBDBDCDCDCDCDCDDDDDDDDDDDDDEDEDEDEDEDFDFDFDFDFDFE0E0E0E0E0),
    .INIT_09(256'hD5D5D5D5D6D6D6D6D6D6D7D7D7D7D7D8D8D8D8D8D9D9D9D9D9D9DADADADADADB),
    .INIT_0A(256'hCFCFCFD0D0D0D0D0D0D1D1D1D1D1D2D2D2D2D2D2D3D3D3D3D3D4D4D4D4D4D4D5),
    .INIT_0B(256'hC9C9C9CACACACACACBCBCBCBCBCBCCCCCCCCCCCDCDCDCDCDCDCECECECECECFCF),
    .INIT_0C(256'hC3C3C4C4C4C4C4C4C5C5C5C5C5C6C6C6C6C6C6C7C7C7C7C7C8C8C8C8C8C9C9C9),
    .INIT_0D(256'hBDBDBEBEBEBEBEBFBFBFBFBFBFC0C0C0C0C0C1C1C1C1C1C2C2C2C2C2C2C3C3C3),
    .INIT_0E(256'hB7B8B8B8B8B8B8B9B9B9B9B9BABABABABABBBBBBBBBBBBBCBCBCBCBCBDBDBDBD),
    .INIT_0F(256'hB1B2B2B2B2B2B3B3B3B3B3B3B4B4B4B4B4B5B5B5B5B5B6B6B6B6B6B6B7B7B7B7),
    .INIT_10(256'hACACACACACACADADADADADAEAEAEAEAEAFAFAFAFAFAFB0B0B0B0B0B1B1B1B1B1),
    .INIT_11(256'hA6A6A6A6A6A7A7A7A7A7A7A8A8A8A8A8A9A9A9A9A9AAAAAAAAAAAAABABABABAB),
    .INIT_12(256'hA0A0A0A0A0A1A1A1A1A1A2A2A2A2A2A2A3A3A3A3A3A4A4A4A4A4A5A5A5A5A5A5),
    .INIT_13(256'h9A9A9A9A9B9B9B9B9B9B9C9C9C9C9C9D9D9D9D9D9D9E9E9E9E9E9F9F9F9F9FA0),
    .INIT_14(256'h949494949595959595959696969696979797979798989898989899999999999A),
    .INIT_15(256'h8E8E8E8E8F8F8F8F8F9090909090909191919191929292929293939393939394),
    .INIT_16(256'h8888888889898989898A8A8A8A8A8B8B8B8B8B8B8C8C8C8C8C8D8D8D8D8D8D8E),
    .INIT_17(256'h8282828383838383838484848484858585858585868686868687878787878888),
    .INIT_18(256'h7C7C7C7D7D7D7D7D7D7E7E7E7E7E7F7F7F7F7F80808080808081818181818282),
    .INIT_19(256'h767676777777777778787878787879797979797A7A7A7A7A7A7B7B7B7B7B7C7C),
    .INIT_1A(256'h7070707171717171727272727272737373737374747474747575757575757676),
    .INIT_1B(256'h6A6A6A6B6B6B6B6B6C6C6C6C6C6C6D6D6D6D6D6E6E6E6E6E6F6F6F6F6F6F7070),
    .INIT_1C(256'h6464646565656565666666666666676767676768686868686969696969696A6A),
    .INIT_1D(256'h5E5E5E5F5F5F5F5F606060606060616161616162626262626363636363636464),
    .INIT_1E(256'h58585859595959595A5A5A5A5A5A5B5B5B5B5B5C5C5C5C5C5D5D5D5D5D5D5E5E),
    .INIT_1F(256'h5252525353535353545454545454555555555556565656565757575757575858),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_012288_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_addra[_o ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i12_008,inst_doa_i12_007,inst_doa_i12_006,inst_doa_i12_005,inst_doa_i12_004,inst_doa_i12_003,inst_doa_i12_002,inst_doa_i12_001,inst_doa_i12_000}));
  // address_offset=13312;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'h4C4C4C4D4D4D4D4D4E4E4E4E4E4E4F4F4F4F4F50505050505151515151515252),
    .INIT_01(256'h464646474747474748484848484849494949494A4A4A4A4A4B4B4B4B4B4B4C4C),
    .INIT_02(256'h4040404141414141414242424242434343434344444444444545454545454646),
    .INIT_03(256'h3A3A3A3B3B3B3B3B3B3C3C3C3C3C3D3D3D3D3D3E3E3E3E3E3E3F3F3F3F3F4040),
    .INIT_04(256'h3434343435353535353636363636373737373738383838383839393939393A3A),
    .INIT_05(256'h2E2E2E2E2F2F2F2F2F3030303030313131313131323232323233333333333434),
    .INIT_06(256'h2828282829292929292A2A2A2A2A2A2B2B2B2B2B2C2C2C2C2C2D2D2D2D2D2E2E),
    .INIT_07(256'h2222222223232323232324242424242525252525262626262627272727272728),
    .INIT_08(256'h1C1C1C1C1C1D1D1D1D1D1E1E1E1E1E1F1F1F1F1F202020202020212121212122),
    .INIT_09(256'h1616161616171717171718181818181919191919191A1A1A1A1A1B1B1B1B1B1C),
    .INIT_0A(256'h1010101010111111111111121212121213131313131414141414151515151515),
    .INIT_0B(256'h0A0A0A0A0A0A0B0B0B0B0B0C0C0C0C0C0D0D0D0D0D0E0E0E0E0E0E0F0F0F0F0F),
    .INIT_0C(256'h0304040404040505050505060606060606070707070708080808080909090909),
    .INIT_0D(256'hFDFEFEFEFEFEFFFFFFFFFFFF0000000000010101010102020202020303030303),
    .INIT_0E(256'hF7F7F8F8F8F8F8F9F9F9F9F9FAFAFAFAFAFBFBFBFBFBFBFCFCFCFCFCFDFDFDFD),
    .INIT_0F(256'hF1F1F2F2F2F2F2F3F3F3F3F3F3F4F4F4F4F4F5F5F5F5F5F6F6F6F6F6F7F7F7F7),
    .INIT_10(256'hEBEBEBECECECECECEDEDEDEDEDEEEEEEEEEEEFEFEFEFEFEFF0F0F0F0F0F1F1F1),
    .INIT_11(256'hE5E5E5E6E6E6E6E6E7E7E7E7E7E7E8E8E8E8E8E9E9E9E9E9EAEAEAEAEAEBEBEB),
    .INIT_12(256'hDFDFDFDFE0E0E0E0E0E1E1E1E1E1E2E2E2E2E2E3E3E3E3E3E3E4E4E4E4E4E5E5),
    .INIT_13(256'hD9D9D9D9DADADADADADBDBDBDBDBDBDCDCDCDCDCDDDDDDDDDDDEDEDEDEDEDFDF),
    .INIT_14(256'hD3D3D3D3D3D4D4D4D4D4D5D5D5D5D5D6D6D6D6D6D6D7D7D7D7D7D8D8D8D8D8D9),
    .INIT_15(256'hCDCDCDCDCDCECECECECECECFCFCFCFCFD0D0D0D0D0D1D1D1D1D1D2D2D2D2D2D2),
    .INIT_16(256'hC6C7C7C7C7C7C8C8C8C8C8C9C9C9C9C9C9CACACACACACBCBCBCBCBCCCCCCCCCC),
    .INIT_17(256'hC0C0C1C1C1C1C1C2C2C2C2C2C3C3C3C3C3C4C4C4C4C4C5C5C5C5C5C5C6C6C6C6),
    .INIT_18(256'hBABABBBBBBBBBBBCBCBCBCBCBCBDBDBDBDBDBEBEBEBEBEBFBFBFBFBFC0C0C0C0),
    .INIT_19(256'hB4B4B4B5B5B5B5B5B6B6B6B6B6B7B7B7B7B7B7B8B8B8B8B8B9B9B9B9B9BABABA),
    .INIT_1A(256'hAEAEAEAEAFAFAFAFAFB0B0B0B0B0B1B1B1B1B1B2B2B2B2B2B3B3B3B3B3B3B4B4),
    .INIT_1B(256'hA8A8A8A8A9A9A9A9A9A9AAAAAAAAAAABABABABABACACACACACADADADADADAEAE),
    .INIT_1C(256'hA2A2A2A2A2A3A3A3A3A3A4A4A4A4A4A4A5A5A5A5A5A6A6A6A6A6A7A7A7A7A7A8),
    .INIT_1D(256'h9B9C9C9C9C9C9D9D9D9D9D9E9E9E9E9E9F9F9F9F9F9FA0A0A0A0A0A1A1A1A1A1),
    .INIT_1E(256'h959596969696969797979797989898989899999999999A9A9A9A9A9A9B9B9B9B),
    .INIT_1F(256'h8F8F909090909090919191919192929292929393939393949494949495959595),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_013312_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_addra[_o ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i13_008,inst_doa_i13_007,inst_doa_i13_006,inst_doa_i13_005,inst_doa_i13_004,inst_doa_i13_003,inst_doa_i13_002,inst_doa_i13_001,inst_doa_i13_000}));
  // address_offset=14336;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'h0000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h8989898A8A8A8A8A8B8B8B8B8B8B8C8C8C8C8C8D8D8D8D8D8E8E8E8E8E8F8F8F),
    .INIT_01(256'h8383838384848484848585858585868686868686878787878788888888888989),
    .INIT_02(256'h7D7D7D7D7D7E7E7E7E7E7F7F7F7F7F8080808080808181818181828282828283),
    .INIT_03(256'h767777777777787878787879797979797A7A7A7A7A7B7B7B7B7B7B7C7C7C7C7C),
    .INIT_04(256'h7070717171717172727272727373737373747474747475757575757676767676),
    .INIT_05(256'h6A6A6A6B6B6B6B6B6C6C6C6C6C6D6D6D6D6D6E6E6E6E6E6F6F6F6F6F70707070),
    .INIT_06(256'h64646465656565656566666666666767676767686868686869696969696A6A6A),
    .INIT_07(256'h5E5E5E5E5F5F5F5F5F5F60606060606161616161626262626263636363636464),
    .INIT_08(256'h58585858585959595959595A5A5A5A5A5B5B5B5B5B5C5C5C5C5C5D5D5D5D5D5E),
    .INIT_09(256'h5152525252525353535353535454545454555555555556565656565757575757),
    .INIT_0A(256'h4B4B4C4C4C4C4C4D4D4D4D4D4D4E4E4E4E4E4F4F4F4F4F505050505051515151),
    .INIT_0B(256'h4545454646464646474747474747484848484849494949494A4A4A4A4A4B4B4B),
    .INIT_0C(256'h3F3F3F3F40404040404041414141414242424242434343434344444444444545),
    .INIT_0D(256'h39393939393A3A3A3A3A3A3B3B3B3B3B3C3C3C3C3C3D3D3D3D3D3E3E3E3E3E3F),
    .INIT_0E(256'h3233333333333434343434343535353535363636363637373737373838383838),
    .INIT_0F(256'h2C2C2D2D2D2D2D2D2E2E2E2E2E2F2F2F2F2F3030303030313131313132323232),
    .INIT_10(256'h262626262727272727282828282829292929292A2A2A2A2A2B2B2B2B2B2C2C2C),
    .INIT_11(256'h2020202020212121212122222222222323232323242424242425252525252626),
    .INIT_12(256'h191A1A1A1A1A1B1B1B1B1B1C1C1C1C1C1D1D1D1D1D1E1E1E1E1E1F1F1F1F1F1F),
    .INIT_13(256'h1313141414141415151515151616161616171717171718181818181819191919),
    .INIT_14(256'h0D0D0D0E0E0E0E0E0F0F0F0F0F10101010101111111111111212121212131313),
    .INIT_15(256'h07070707080808080809090909090A0A0A0A0A0A0B0B0B0B0B0C0C0C0C0C0D0D),
    .INIT_16(256'h0101010101020202020203030303030304040404040505050505060606060607),
    .INIT_17(256'hFAFBFBFBFBFBFBFCFCFCFCFCFDFDFDFDFDFEFEFEFEFEFFFFFFFFFF0000000000),
    .INIT_18(256'hF4F4F4F5F5F5F5F5F6F6F6F6F6F7F7F7F7F7F8F8F8F8F8F9F9F9F9F9FAFAFAFA),
    .INIT_19(256'hEEEEEEEEEFEFEFEFEFF0F0F0F0F0F1F1F1F1F1F2F2F2F2F2F3F3F3F3F3F4F4F4),
    .INIT_1A(256'hE8E8E8E8E8E9E9E9E9E9EAEAEAEAEAEBEBEBEBEBECECECECECECEDEDEDEDEDEE),
    .INIT_1B(256'hE1E2E2E2E2E2E3E3E3E3E3E4E4E4E4E4E4E5E5E5E5E5E6E6E6E6E6E7E7E7E7E7),
    .INIT_1C(256'hDBDBDCDCDCDCDCDCDDDDDDDDDDDEDEDEDEDEDFDFDFDFDFE0E0E0E0E0E1E1E1E1),
    .INIT_1D(256'hD5D5D5D5D6D6D6D6D6D7D7D7D7D7D8D8D8D8D8D9D9D9D9D9DADADADADADBDBDB),
    .INIT_1E(256'hCFCFCFCFCFD0D0D0D0D0D1D1D1D1D1D2D2D2D2D2D3D3D3D3D3D4D4D4D4D4D4D5),
    .INIT_1F(256'hC8C9C9C9C9C9CACACACACACBCBCBCBCBCCCCCCCCCCCCCDCDCDCDCDCECECECECE),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_014336_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_addra[_o ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i14_008,inst_doa_i14_007,inst_doa_i14_006,inst_doa_i14_005,inst_doa_i14_004,inst_doa_i14_003,inst_doa_i14_002,inst_doa_i14_001,inst_doa_i14_000}));
  // address_offset=15360;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hC2C2C3C3C3C3C3C4C4C4C4C4C4C5C5C5C5C5C6C6C6C6C6C7C7C7C7C7C8C8C8C8),
    .INIT_01(256'hBCBCBCBCBDBDBDBDBDBEBEBEBEBEBFBFBFBFBFC0C0C0C0C0C1C1C1C1C1C2C2C2),
    .INIT_02(256'hB6B6B6B6B6B7B7B7B7B7B8B8B8B8B8B9B9B9B9B9BABABABABABBBBBBBBBBBBBC),
    .INIT_03(256'hAFB0B0B0B0B0B1B1B1B1B1B2B2B2B2B2B2B3B3B3B3B3B4B4B4B4B4B5B5B5B5B5),
    .INIT_04(256'hA9A9A9AAAAAAAAAAABABABABABACACACACACADADADADADAEAEAEAEAEAFAFAFAF),
    .INIT_05(256'hA3A3A3A3A4A4A4A4A4A5A5A5A5A5A6A6A6A6A6A7A7A7A7A7A8A8A8A8A8A9A9A9),
    .INIT_06(256'h9D9D9D9D9D9E9E9E9E9E9F9F9F9F9FA0A0A0A0A0A0A1A1A1A1A1A2A2A2A2A2A3),
    .INIT_07(256'h96979797979797989898989899999999999A9A9A9A9A9B9B9B9B9B9C9C9C9C9C),
    .INIT_08(256'h9090909191919191929292929293939393939494949494959595959596969696),
    .INIT_09(256'h8A8A8A8A8B8B8B8B8B8C8C8C8C8C8D8D8D8D8D8E8E8E8E8E8E8F8F8F8F8F9090),
    .INIT_0A(256'h848484848484858585858586868686868787878787888888888889898989898A),
    .INIT_0B(256'h7D7D7E7E7E7E7E7F7F7F7F7F8080808080818181818182828282828383838383),
    .INIT_0C(256'h777777787878787879797979797A7A7A7A7A7B7B7B7B7B7B7C7C7C7C7C7D7D7D),
    .INIT_0D(256'h7171717171727272727273737373737474747474757575757576767676767777),
    .INIT_0E(256'h6A6B6B6B6B6B6C6C6C6C6C6D6D6D6D6D6E6E6E6E6E6F6F6F6F6F707070707071),
    .INIT_0F(256'h646465656565656666666666676767676767686868686869696969696A6A6A6A),
    .INIT_10(256'h5E5E5E5E5F5F5F5F5F6060606060616161616162626262626363636363646464),
    .INIT_11(256'h585858585859595959595A5A5A5A5A5B5B5B5B5B5C5C5C5C5C5D5D5D5D5D5D5E),
    .INIT_12(256'h5152525252525353535353535454545454555555555556565656565757575757),
    .INIT_13(256'h4B4B4B4C4C4C4C4C4D4D4D4D4D4E4E4E4E4E4F4F4F4F4F505050505051515151),
    .INIT_14(256'h454545454646464646474747474748484848484949494949494A4A4A4A4A4B4B),
    .INIT_15(256'h3F3F3F3F3F3F4040404040414141414142424242424343434343444444444445),
    .INIT_16(256'h383839393939393A3A3A3A3A3B3B3B3B3B3C3C3C3C3C3D3D3D3D3D3E3E3E3E3E),
    .INIT_17(256'h3232323333333333343434343434353535353536363636363737373737383838),
    .INIT_18(256'h2C2C2C2C2C2D2D2D2D2D2E2E2E2E2E2F2F2F2F2F303030303031313131313232),
    .INIT_19(256'h2526262626262727272727282828282829292929292A2A2A2A2A2A2B2B2B2B2B),
    .INIT_1A(256'h1F1F1F2020202020212121212122222222222323232323242424242425252525),
    .INIT_1B(256'h191919191A1A1A1A1A1B1B1B1B1B1C1C1C1C1C1D1D1D1D1D1E1E1E1E1E1F1F1F),
    .INIT_1C(256'h1313131313141414141415151515151516161616161717171717181818181819),
    .INIT_1D(256'h0C0C0D0D0D0D0D0E0E0E0E0E0F0F0F0F0F101010101011111111111212121212),
    .INIT_1E(256'h0606060707070707080808080809090909090A0A0A0A0A0A0B0B0B0B0B0C0C0C),
    .INIT_1F(256'h0000000000010101010102020202020303030303040404040405050505050606),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_015360_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_addra[_o ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i15_008,inst_doa_i15_007,inst_doa_i15_006,inst_doa_i15_005,inst_doa_i15_004,inst_doa_i15_003,inst_doa_i15_002,inst_doa_i15_001,inst_doa_i15_000}));
  // address_offset=16384;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'hF9FAFAFAFAFAFBFBFBFBFBFCFCFCFCFCFDFDFDFDFDFEFEFEFEFEFFFFFFFFFFFF),
    .INIT_01(256'hF3F3F4F4F4F4F4F5F5F5F5F5F5F6F6F6F6F6F7F7F7F7F7F8F8F8F8F8F9F9F9F9),
    .INIT_02(256'hEDEDEDEDEEEEEEEEEEEFEFEFEFEFF0F0F0F0F0F1F1F1F1F1F2F2F2F2F2F3F3F3),
    .INIT_03(256'hE7E7E7E7E7E8E8E8E8E8E9E9E9E9E9EAEAEAEAEAEAEBEBEBEBEBECECECECECED),
    .INIT_04(256'hE0E0E1E1E1E1E1E2E2E2E2E2E3E3E3E3E3E4E4E4E4E4E5E5E5E5E5E6E6E6E6E6),
    .INIT_05(256'hDADADADBDBDBDBDBDCDCDCDCDCDDDDDDDDDDDEDEDEDEDEDFDFDFDFDFE0E0E0E0),
    .INIT_06(256'hD4D4D4D4D5D5D5D5D5D5D6D6D6D6D6D7D7D7D7D7D8D8D8D8D8D9D9D9D9D9DADA),
    .INIT_07(256'hCDCECECECECECFCFCFCFCFD0D0D0D0D0D1D1D1D1D1D2D2D2D2D2D3D3D3D3D3D4),
    .INIT_08(256'hC7C7C8C8C8C8C8C9C9C9C9C9CACACACACACBCBCBCBCBCBCCCCCCCCCCCDCDCDCD),
    .INIT_09(256'hC1C1C1C1C2C2C2C2C2C3C3C3C3C3C4C4C4C4C4C5C5C5C5C5C6C6C6C6C6C7C7C7),
    .INIT_0A(256'hBBBBBBBBBBBCBCBCBCBCBDBDBDBDBDBEBEBEBEBEBFBFBFBFBFC0C0C0C0C0C0C1),
    .INIT_0B(256'hB4B5B5B5B5B5B6B6B6B6B6B6B7B7B7B7B7B8B8B8B8B8B9B9B9B9B9BABABABABA),
    .INIT_0C(256'hAEAEAEAFAFAFAFAFB0B0B0B0B0B1B1B1B1B1B2B2B2B2B2B3B3B3B3B3B4B4B4B4),
    .INIT_0D(256'hA8A8A8A8A9A9A9A9A9AAAAAAAAAAABABABABABACACACACACACADADADADADAEAE),
    .INIT_0E(256'hA2A2A2A2A2A2A3A3A3A3A3A4A4A4A4A4A5A5A5A5A5A6A6A6A6A6A7A7A7A7A7A8),
    .INIT_0F(256'h9B9B9C9C9C9C9C9D9D9D9D9D9E9E9E9E9E9F9F9F9F9FA0A0A0A0A0A1A1A1A1A1),
    .INIT_10(256'h9595959696969696979797979798989898989899999999999A9A9A9A9A9B9B9B),
    .INIT_11(256'h8F8F8F8F8F909090909091919191919292929292939393939394949494949595),
    .INIT_12(256'h8889898989898A8A8A8A8A8B8B8B8B8B8C8C8C8C8C8D8D8D8D8D8E8E8E8E8E8E),
    .INIT_13(256'h8282838383838384848484848485858585858686868686878787878788888888),
    .INIT_14(256'h7C7C7C7C7D7D7D7D7D7E7E7E7E7E7F7F7F7F7F80808080808181818181828282),
    .INIT_15(256'h76767676767777777777787878787879797979797A7A7A7A7A7B7B7B7B7B7B7C),
    .INIT_16(256'h6F70707070707171717171717272727272737373737374747474747575757575),
    .INIT_17(256'h6969696A6A6A6A6A6B6B6B6B6B6C6C6C6C6C6D6D6D6D6D6E6E6E6E6E6F6F6F6F),
    .INIT_18(256'h6363636364646464646565656565666666666667676767676868686868686969),
    .INIT_19(256'h5D5D5D5D5D5E5E5E5E5E5F5F5F5F5F5F60606060606161616161626262626263),
    .INIT_1A(256'h56565757575757585858585859595959595A5A5A5A5A5B5B5B5B5B5C5C5C5C5C),
    .INIT_1B(256'h5050505151515151525252525253535353535454545454555555555556565656),
    .INIT_1C(256'h4A4A4A4A4B4B4B4B4B4C4C4C4C4C4D4D4D4D4D4D4E4E4E4E4E4F4F4F4F4F5050),
    .INIT_1D(256'h444444444444454545454546464646464747474747484848484849494949494A),
    .INIT_1E(256'h3D3D3E3E3E3E3E3F3F3F3F3F4040404040414141414142424242424343434343),
    .INIT_1F(256'h373737383838383839393939393A3A3A3A3A3B3B3B3B3B3B3C3C3C3C3C3D3D3D),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_016384_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_Naddr_o_al_n28 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i16_008,inst_doa_i16_007,inst_doa_i16_006,inst_doa_i16_005,inst_doa_i16_004,inst_doa_i16_003,inst_doa_i16_002,inst_doa_i16_001,inst_doa_i16_000}));
  // address_offset=16384;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'h000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_016384_009 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n1070,open_n1071,open_n1072,open_n1073,open_n1074,open_n1075,open_n1076,1'b0,open_n1077}),
    .rsta(rsta),
    .doa({open_n1092,open_n1093,open_n1094,open_n1095,open_n1096,open_n1097,open_n1098,open_n1099,inst_doa_i16_009}));
  // address_offset=16384;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'h0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_016384_010 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n1128,open_n1129,open_n1130,open_n1131,open_n1132,open_n1133,open_n1134,1'b0,open_n1135}),
    .rsta(rsta),
    .doa({open_n1150,open_n1151,open_n1152,open_n1153,open_n1154,open_n1155,open_n1156,open_n1157,inst_doa_i16_010}));
  // address_offset=16384;data_offset=11;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_016384_011 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n1186,open_n1187,open_n1188,open_n1189,open_n1190,open_n1191,open_n1192,1'b0,open_n1193}),
    .rsta(rsta),
    .doa({open_n1208,open_n1209,open_n1210,open_n1211,open_n1212,open_n1213,open_n1214,open_n1215,inst_doa_i16_011}));
  // address_offset=17408;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'h000000000000000000000000000000000000000000000000000000000FFFFFFF),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h3131313132323232323333333333333434343434353535353536363636363737),
    .INIT_01(256'h2B2B2B2B2B2B2C2C2C2C2C2D2D2D2D2D2E2E2E2E2E2F2F2F2F2F303030303031),
    .INIT_02(256'h2424252525252526262626262727272727282828282829292929292A2A2A2A2A),
    .INIT_03(256'h1E1E1E1F1F1F1F1F202020202021212121212222222222232323232323242424),
    .INIT_04(256'h1818181819191919191A1A1A1A1A1B1B1B1B1B1B1C1C1C1C1C1D1D1D1D1D1E1E),
    .INIT_05(256'h1212121212131313131313141414141415151515151616161616171717171718),
    .INIT_06(256'h0B0B0C0C0C0C0C0D0D0D0D0D0E0E0E0E0E0F0F0F0F0F10101010101111111111),
    .INIT_07(256'h05050506060606060707070707080808080809090909090A0A0A0A0A0B0B0B0B),
    .INIT_08(256'hFFFFFFFF00000000000101010101020202020203030303030404040404040505),
    .INIT_09(256'hF9F9F9F9F9FAFAFAFAFAFBFBFBFBFBFCFCFCFCFCFCFDFDFDFDFDFEFEFEFEFEFF),
    .INIT_0A(256'hF2F3F3F3F3F3F4F4F4F4F4F5F5F5F5F5F5F6F6F6F6F6F7F7F7F7F7F8F8F8F8F8),
    .INIT_0B(256'hECECEDEDEDEDEDEEEEEEEEEEEEEFEFEFEFEFF0F0F0F0F0F1F1F1F1F1F2F2F2F2),
    .INIT_0C(256'hE6E6E6E7E7E7E7E7E7E8E8E8E8E8E9E9E9E9E9EAEAEAEAEAEBEBEBEBEBECECEC),
    .INIT_0D(256'hE0E0E0E0E0E1E1E1E1E1E2E2E2E2E2E3E3E3E3E3E4E4E4E4E4E5E5E5E5E5E6E6),
    .INIT_0E(256'hD9DADADADADADBDBDBDBDBDCDCDCDCDCDDDDDDDDDDDEDEDEDEDEDFDFDFDFDFE0),
    .INIT_0F(256'hD3D3D4D4D4D4D4D5D5D5D5D5D6D6D6D6D6D7D7D7D7D7D8D8D8D8D8D9D9D9D9D9),
    .INIT_10(256'hCDCDCDCECECECECECFCFCFCFCFD0D0D0D0D0D1D1D1D1D1D2D2D2D2D2D2D3D3D3),
    .INIT_11(256'hC7C7C7C7C8C8C8C8C8C9C9C9C9C9CACACACACACBCBCBCBCBCBCCCCCCCCCCCDCD),
    .INIT_12(256'hC1C1C1C1C1C2C2C2C2C2C3C3C3C3C3C4C4C4C4C4C5C5C5C5C5C5C6C6C6C6C6C7),
    .INIT_13(256'hBABBBBBBBBBBBCBCBCBCBCBDBDBDBDBDBEBEBEBEBEBFBFBFBFBFBFC0C0C0C0C0),
    .INIT_14(256'hB4B4B5B5B5B5B5B6B6B6B6B6B7B7B7B7B7B8B8B8B8B8B8B9B9B9B9B9BABABABA),
    .INIT_15(256'hAEAEAEAFAFAFAFAFB0B0B0B0B0B1B1B1B1B1B2B2B2B2B2B2B3B3B3B3B3B4B4B4),
    .INIT_16(256'hA8A8A8A8A9A9A9A9A9AAAAAAAAAAABABABABABACACACACACACADADADADADAEAE),
    .INIT_17(256'hA2A2A2A2A2A3A3A3A3A3A4A4A4A4A4A5A5A5A5A5A6A6A6A6A6A6A7A7A7A7A7A8),
    .INIT_18(256'h9B9C9C9C9C9C9D9D9D9D9D9E9E9E9E9E9F9F9F9F9FA0A0A0A0A0A0A1A1A1A1A1),
    .INIT_19(256'h959596969696969797979797989898989899999999999A9A9A9A9A9A9B9B9B9B),
    .INIT_1A(256'h8F8F8F9090909090919191919192929292929393939393949494949495959595),
    .INIT_1B(256'h898989898A8A8A8A8A8B8B8B8B8B8C8C8C8C8C8D8D8D8D8D8E8E8E8E8E8F8F8F),
    .INIT_1C(256'h8383838384848484848485858585858686868686878787878788888888888989),
    .INIT_1D(256'h7D7D7D7D7D7E7E7E7E7E7F7F7F7F7F7F80808080808181818181828282828283),
    .INIT_1E(256'h76777777777778787878787979797979797A7A7A7A7A7B7B7B7B7B7C7C7C7C7C),
    .INIT_1F(256'h7070717171717172727272727373737373747474747474757575757576767676),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_017408_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_Naddr_o_al_n28 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i17_008,inst_doa_i17_007,inst_doa_i17_006,inst_doa_i17_005,inst_doa_i17_004,inst_doa_i17_003,inst_doa_i17_002,inst_doa_i17_001,inst_doa_i17_000}));
  // address_offset=18432;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'h6A6A6A6B6B6B6B6B6C6C6C6C6C6D6D6D6D6D6E6E6E6E6E6F6F6F6F6F6F707070),
    .INIT_01(256'h64646465656565656566666666666767676767686868686869696969696A6A6A),
    .INIT_02(256'h5E5E5E5E5F5F5F5F5F6060606060606161616161626262626263636363636464),
    .INIT_03(256'h585858585859595959595A5A5A5A5A5B5B5B5B5B5B5C5C5C5C5C5D5D5D5D5D5E),
    .INIT_04(256'h5152525252525353535353545454545455555555555656565656565757575757),
    .INIT_05(256'h4B4C4C4C4C4C4C4D4D4D4D4D4E4E4E4E4E4F4F4F4F4F50505050505151515151),
    .INIT_06(256'h45454646464646474747474748484848484849494949494A4A4A4A4A4B4B4B4B),
    .INIT_07(256'h3F3F3F4040404040414141414142424242424343434343434444444444454545),
    .INIT_08(256'h3939393A3A3A3A3A3A3B3B3B3B3B3C3C3C3C3C3D3D3D3D3D3E3E3E3E3E3F3F3F),
    .INIT_09(256'h3333333334343434343535353535363636363636373737373738383838383939),
    .INIT_0A(256'h2D2D2D2D2D2E2E2E2E2E2F2F2F2F2F3030303030313131313131323232323233),
    .INIT_0B(256'h272727272728282828282929292929292A2A2A2A2A2B2B2B2B2B2C2C2C2C2C2D),
    .INIT_0C(256'h2021212121212222222222232323232324242424242425252525252626262626),
    .INIT_0D(256'h1A1B1B1B1B1B1C1C1C1C1C1C1D1D1D1D1D1E1E1E1E1E1F1F1F1F1F2020202020),
    .INIT_0E(256'h141415151515151616161616171717171718181818181819191919191A1A1A1A),
    .INIT_0F(256'h0E0E0F0F0F0F0F10101010101011111111111212121212131313131314141414),
    .INIT_10(256'h08080809090909090A0A0A0A0A0B0B0B0B0B0C0C0C0C0C0C0D0D0D0D0D0E0E0E),
    .INIT_11(256'h0202020303030303040404040404050505050506060606060707070707080808),
    .INIT_12(256'hFCFCFCFCFDFDFDFDFDFEFEFEFEFEFFFFFFFFFF00000000000001010101010202),
    .INIT_13(256'hF6F6F6F6F7F7F7F7F7F8F8F8F8F8F9F9F9F9F9F9FAFAFAFAFAFBFBFBFBFBFCFC),
    .INIT_14(256'hF0F0F0F0F1F1F1F1F1F1F2F2F2F2F2F3F3F3F3F3F4F4F4F4F4F5F5F5F5F5F5F6),
    .INIT_15(256'hEAEAEAEAEAEBEBEBEBEBECECECECECEDEDEDEDEDEEEEEEEEEEEEEFEFEFEFEFF0),
    .INIT_16(256'hE4E4E4E4E4E5E5E5E5E5E6E6E6E6E6E6E7E7E7E7E7E8E8E8E8E8E9E9E9E9E9EA),
    .INIT_17(256'hDEDEDEDEDEDFDFDFDFDFDFE0E0E0E0E0E1E1E1E1E1E2E2E2E2E2E3E3E3E3E3E3),
    .INIT_18(256'hD8D8D8D8D8D8D9D9D9D9D9DADADADADADBDBDBDBDBDCDCDCDCDCDCDDDDDDDDDD),
    .INIT_19(256'hD1D2D2D2D2D2D3D3D3D3D3D4D4D4D4D4D5D5D5D5D5D5D6D6D6D6D6D7D7D7D7D7),
    .INIT_1A(256'hCBCCCCCCCCCCCDCDCDCDCDCECECECECECECFCFCFCFCFD0D0D0D0D0D1D1D1D1D1),
    .INIT_1B(256'hC5C6C6C6C6C6C7C7C7C7C7C7C8C8C8C8C8C9C9C9C9C9CACACACACACBCBCBCBCB),
    .INIT_1C(256'hBFC0C0C0C0C0C1C1C1C1C1C1C2C2C2C2C2C3C3C3C3C3C4C4C4C4C4C4C5C5C5C5),
    .INIT_1D(256'hB9BABABABABABABBBBBBBBBBBCBCBCBCBCBDBDBDBDBDBEBEBEBEBEBEBFBFBFBF),
    .INIT_1E(256'hB3B4B4B4B4B4B4B5B5B5B5B5B6B6B6B6B6B7B7B7B7B7B7B8B8B8B8B8B9B9B9B9),
    .INIT_1F(256'hADAEAEAEAEAEAEAFAFAFAFAFB0B0B0B0B0B1B1B1B1B1B1B2B2B2B2B2B3B3B3B3),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_018432_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_Naddr_o_al_n28 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i18_008,inst_doa_i18_007,inst_doa_i18_006,inst_doa_i18_005,inst_doa_i18_004,inst_doa_i18_003,inst_doa_i18_002,inst_doa_i18_001,inst_doa_i18_000}));
  // address_offset=19456;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'h0000000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'hA7A8A8A8A8A8A8A9A9A9A9A9AAAAAAAAAAABABABABABABACACACACACADADADAD),
    .INIT_01(256'hA1A2A2A2A2A2A2A3A3A3A3A3A4A4A4A4A4A5A5A5A5A5A5A6A6A6A6A6A7A7A7A7),
    .INIT_02(256'h9B9C9C9C9C9C9C9D9D9D9D9D9E9E9E9E9E9F9F9F9F9F9FA0A0A0A0A0A1A1A1A1),
    .INIT_03(256'h95969696969696979797979798989898989999999999999A9A9A9A9A9B9B9B9B),
    .INIT_04(256'h8F90909090909091919191919292929292939393939393949494949495959595),
    .INIT_05(256'h898A8A8A8A8A8A8B8B8B8B8B8C8C8C8C8C8D8D8D8D8D8D8E8E8E8E8E8F8F8F8F),
    .INIT_06(256'h8384848484848585858585858686868686878787878787888888888889898989),
    .INIT_07(256'h7D7E7E7E7E7E7F7F7F7F7F7F8080808080818181818182828282828283838383),
    .INIT_08(256'h77787878787879797979797A7A7A7A7A7A7B7B7B7B7B7C7C7C7C7C7C7D7D7D7D),
    .INIT_09(256'h7272727272727373737373747474747474757575757576767676767777777777),
    .INIT_0A(256'h6C6C6C6C6C6C6D6D6D6D6D6E6E6E6E6E6F6F6F6F6F6F70707070707171717171),
    .INIT_0B(256'h6666666666676767676767686868686869696969696A6A6A6A6A6A6B6B6B6B6B),
    .INIT_0C(256'h6060606060616161616162626262626263636363636464646464646565656565),
    .INIT_0D(256'h5A5A5A5A5A5B5B5B5B5B5C5C5C5C5C5D5D5D5D5D5D5E5E5E5E5E5F5F5F5F5F5F),
    .INIT_0E(256'h545454545555555555555656565656575757575758585858585859595959595A),
    .INIT_0F(256'h4E4E4E4E4F4F4F4F4F5050505050505151515151525252525253535353535354),
    .INIT_10(256'h4848484949494949494A4A4A4A4A4B4B4B4B4B4C4C4C4C4C4C4D4D4D4D4D4E4E),
    .INIT_11(256'h4242424343434343444444444444454545454546464646464747474747474848),
    .INIT_12(256'h3C3C3D3D3D3D3D3D3E3E3E3E3E3F3F3F3F3F4040404040404141414141424242),
    .INIT_13(256'h3636373737373738383838383939393939393A3A3A3A3A3B3B3B3B3B3B3C3C3C),
    .INIT_14(256'h3031313131313232323232323333333333343434343434353535353536363636),
    .INIT_15(256'h2B2B2B2B2B2B2C2C2C2C2C2D2D2D2D2D2D2E2E2E2E2E2F2F2F2F2F2F30303030),
    .INIT_16(256'h2525252525262626262626272727272728282828282929292929292A2A2A2A2A),
    .INIT_17(256'h1F1F1F1F20202020202021212121212222222222222323232323242424242424),
    .INIT_18(256'h191919191A1A1A1A1A1B1B1B1B1B1C1C1C1C1C1C1D1D1D1D1D1E1E1E1E1E1E1F),
    .INIT_19(256'h1313131414141414151515151515161616161617171717171718181818181919),
    .INIT_1A(256'h0D0D0E0E0E0E0E0F0F0F0F0F0F10101010101111111111111212121212131313),
    .INIT_1B(256'h0708080808080909090909090A0A0A0A0A0B0B0B0B0B0B0C0C0C0C0C0D0D0D0D),
    .INIT_1C(256'h0202020202020303030303040404040404050505050506060606060607070707),
    .INIT_1D(256'hFCFCFCFCFCFDFDFDFDFDFEFEFEFEFEFEFFFFFFFFFF0000000000000101010101),
    .INIT_1E(256'hF6F6F6F6F7F7F7F7F7F8F8F8F8F8F8F9F9F9F9F9FAFAFAFAFAFAFBFBFBFBFBFC),
    .INIT_1F(256'hF0F0F0F1F1F1F1F1F2F2F2F2F2F2F3F3F3F3F3F4F4F4F4F4F4F5F5F5F5F5F6F6),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_019456_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_Naddr_o_al_n28 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i19_008,inst_doa_i19_007,inst_doa_i19_006,inst_doa_i19_005,inst_doa_i19_004,inst_doa_i19_003,inst_doa_i19_002,inst_doa_i19_001,inst_doa_i19_000}));
  // address_offset=20480;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hEAEBEBEBEBEBEBECECECECECEDEDEDEDEDEDEEEEEEEEEEEFEFEFEFEFEFF0F0F0),
    .INIT_01(256'hE5E5E5E5E5E5E6E6E6E6E6E7E7E7E7E7E7E8E8E8E8E8E9E9E9E9E9E9EAEAEAEA),
    .INIT_02(256'hDFDFDFDFDFE0E0E0E0E0E1E1E1E1E1E1E2E2E2E2E2E3E3E3E3E3E3E4E4E4E4E4),
    .INIT_03(256'hD9D9D9DADADADADADADBDBDBDBDBDCDCDCDCDCDCDDDDDDDDDDDDDEDEDEDEDEDF),
    .INIT_04(256'hD3D3D4D4D4D4D4D4D5D5D5D5D5D6D6D6D6D6D6D7D7D7D7D7D8D8D8D8D8D8D9D9),
    .INIT_05(256'hCDCECECECECECFCFCFCFCFCFD0D0D0D0D0D1D1D1D1D1D1D2D2D2D2D2D2D3D3D3),
    .INIT_06(256'hC8C8C8C8C8C9C9C9C9C9C9CACACACACACBCBCBCBCBCBCCCCCCCCCCCDCDCDCDCD),
    .INIT_07(256'hC2C2C2C2C3C3C3C3C3C4C4C4C4C4C4C5C5C5C5C5C6C6C6C6C6C6C7C7C7C7C7C8),
    .INIT_08(256'hBCBCBDBDBDBDBDBDBEBEBEBEBEBFBFBFBFBFBFC0C0C0C0C0C1C1C1C1C1C1C2C2),
    .INIT_09(256'hB6B7B7B7B7B7B8B8B8B8B8B8B9B9B9B9B9BABABABABABABBBBBBBBBBBBBCBCBC),
    .INIT_0A(256'hB1B1B1B1B1B2B2B2B2B2B3B3B3B3B3B3B4B4B4B4B4B5B5B5B5B5B5B6B6B6B6B6),
    .INIT_0B(256'hABABABACACACACACACADADADADADAEAEAEAEAEAEAFAFAFAFAFB0B0B0B0B0B0B1),
    .INIT_0C(256'hA5A6A6A6A6A6A6A7A7A7A7A7A7A8A8A8A8A8A9A9A9A9A9A9AAAAAAAAAAABABAB),
    .INIT_0D(256'hA0A0A0A0A0A1A1A1A1A1A1A2A2A2A2A2A2A3A3A3A3A3A4A4A4A4A4A4A5A5A5A5),
    .INIT_0E(256'h9A9A9A9A9B9B9B9B9B9C9C9C9C9C9C9D9D9D9D9D9D9E9E9E9E9E9F9F9F9F9F9F),
    .INIT_0F(256'h9494959595959596969696969697979797979798989898989999999999999A9A),
    .INIT_10(256'h8F8F8F8F8F8F9090909090919191919191929292929292939393939394949494),
    .INIT_11(256'h898989898A8A8A8A8A8B8B8B8B8B8B8C8C8C8C8C8C8D8D8D8D8D8E8E8E8E8E8E),
    .INIT_12(256'h8383848484848484858585858586868686868687878787878888888888888989),
    .INIT_13(256'h7E7E7E7E7E7E7F7F7F7F7F808080808080818181818181828282828283838383),
    .INIT_14(256'h7878787879797979797A7A7A7A7A7A7B7B7B7B7B7B7C7C7C7C7C7D7D7D7D7D7D),
    .INIT_15(256'h7273737373737374747474747475757575757676767676767777777777777878),
    .INIT_16(256'h6D6D6D6D6D6E6E6E6E6E6E6F6F6F6F6F70707070707071717171717172727272),
    .INIT_17(256'h67676768686868686869696969696A6A6A6A6A6A6B6B6B6B6B6B6C6C6C6C6C6D),
    .INIT_18(256'h6162626262626363636363636464646464646565656565666666666666676767),
    .INIT_19(256'h5C5C5C5C5D5D5D5D5D5D5E5E5E5E5E5F5F5F5F5F5F6060606060606161616161),
    .INIT_1A(256'h565657575757575858585858585959595959595A5A5A5A5A5A5B5B5B5B5B5C5C),
    .INIT_1B(256'h5151515151525252525252535353535354545454545455555555555556565656),
    .INIT_1C(256'h4B4B4B4C4C4C4C4C4D4D4D4D4D4D4E4E4E4E4E4E4F4F4F4F4F50505050505051),
    .INIT_1D(256'h46464646464647474747474748484848484949494949494A4A4A4A4A4A4B4B4B),
    .INIT_1E(256'h4040404141414141414242424242424343434343444444444444454545454545),
    .INIT_1F(256'h3A3B3B3B3B3B3C3C3C3C3C3C3D3D3D3D3D3D3E3E3E3E3E3E3F3F3F3F3F404040),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_020480_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_Naddra_o_al_n36 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i20_008,inst_doa_i20_007,inst_doa_i20_006,inst_doa_i20_005,inst_doa_i20_004,inst_doa_i20_003,inst_doa_i20_002,inst_doa_i20_001,inst_doa_i20_000}));
  // address_offset=21504;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'h3535353536363636363737373737373838383838383939393939393A3A3A3A3A),
    .INIT_01(256'h2F30303030303031313131313132323232323333333333333434343434343535),
    .INIT_02(256'h2A2A2A2A2B2B2B2B2B2B2C2C2C2C2C2C2D2D2D2D2D2E2E2E2E2E2E2F2F2F2F2F),
    .INIT_03(256'h2425252525252526262626262627272727272728282828282929292929292A2A),
    .INIT_04(256'h1F1F1F1F20202020202021212121212122222222222323232323232424242424),
    .INIT_05(256'h191A1A1A1A1A1A1B1B1B1B1B1B1C1C1C1C1C1C1D1D1D1D1D1E1E1E1E1E1E1F1F),
    .INIT_06(256'h1414141415151515151516161616161617171717171818181818181919191919),
    .INIT_07(256'h0E0F0F0F0F0F0F10101010101111111111111212121212121313131313131414),
    .INIT_08(256'h0909090A0A0A0A0A0A0B0B0B0B0B0B0C0C0C0C0C0C0D0D0D0D0D0D0E0E0E0E0E),
    .INIT_09(256'h0404040404040505050505050606060606060707070707070808080808080909),
    .INIT_0A(256'hFEFEFEFFFFFFFFFFFF0000000000000101010101020202020202030303030303),
    .INIT_0B(256'hF9F9F9F9F9FAFAFAFAFAFAFBFBFBFBFBFBFCFCFCFCFCFCFDFDFDFDFDFDFEFEFE),
    .INIT_0C(256'hF3F3F4F4F4F4F4F4F5F5F5F5F5F5F6F6F6F6F6F6F7F7F7F7F7F7F8F8F8F8F8F9),
    .INIT_0D(256'hEEEEEEEEEFEFEFEFEFEFF0F0F0F0F0F0F1F1F1F1F1F1F2F2F2F2F2F2F3F3F3F3),
    .INIT_0E(256'hE8E9E9E9E9E9E9EAEAEAEAEAEAEBEBEBEBEBEBECECECECECECEDEDEDEDEDEEEE),
    .INIT_0F(256'hE3E3E3E4E4E4E4E4E4E5E5E5E5E5E5E6E6E6E6E6E6E7E7E7E7E7E7E8E8E8E8E8),
    .INIT_10(256'hDEDEDEDEDEDFDFDFDFDFDFE0E0E0E0E0E0E1E1E1E1E1E1E2E2E2E2E2E2E3E3E3),
    .INIT_11(256'hD8D8D9D9D9D9D9D9DADADADADADADBDBDBDBDBDBDCDCDCDCDCDCDDDDDDDDDDDD),
    .INIT_12(256'hD3D3D3D3D4D4D4D4D4D4D5D5D5D5D5D5D6D6D6D6D6D6D7D7D7D7D7D7D8D8D8D8),
    .INIT_13(256'hCECECECECECECFCFCFCFCFCFD0D0D0D0D0D0D1D1D1D1D1D1D2D2D2D2D2D2D3D3),
    .INIT_14(256'hC8C8C9C9C9C9C9C9CACACACACACACBCBCBCBCBCBCCCCCCCCCCCCCDCDCDCDCDCD),
    .INIT_15(256'hC3C3C3C3C4C4C4C4C4C4C5C5C5C5C5C5C6C6C6C6C6C6C7C7C7C7C7C7C8C8C8C8),
    .INIT_16(256'hBEBEBEBEBEBEBFBFBFBFBFBFC0C0C0C0C0C0C1C1C1C1C1C1C2C2C2C2C2C2C3C3),
    .INIT_17(256'hB8B8B9B9B9B9B9B9BABABABABABABBBBBBBBBBBBBCBCBCBCBCBCBDBDBDBDBDBD),
    .INIT_18(256'hB3B3B3B3B4B4B4B4B4B4B5B5B5B5B5B5B6B6B6B6B6B6B7B7B7B7B7B7B8B8B8B8),
    .INIT_19(256'hAEAEAEAEAEAEAFAFAFAFAFAFB0B0B0B0B0B0B1B1B1B1B1B1B2B2B2B2B2B2B3B3),
    .INIT_1A(256'hA8A9A9A9A9A9A9AAAAAAAAAAAAABABABABABABACACACACACACADADADADADADAD),
    .INIT_1B(256'hA3A3A3A4A4A4A4A4A4A5A5A5A5A5A5A6A6A6A6A6A6A7A7A7A7A7A7A8A8A8A8A8),
    .INIT_1C(256'h9E9E9E9E9F9F9F9F9F9F9FA0A0A0A0A0A0A1A1A1A1A1A1A2A2A2A2A2A2A3A3A3),
    .INIT_1D(256'h9999999999999A9A9A9A9A9A9B9B9B9B9B9B9C9C9C9C9C9C9D9D9D9D9D9D9E9E),
    .INIT_1E(256'h9394949494949495959595959595969696969696979797979797989898989898),
    .INIT_1F(256'h8E8E8E8F8F8F8F8F8F9090909090909191919191919292929292929393939393),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_021504_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_Naddra_o_al_n36 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i21_008,inst_doa_i21_007,inst_doa_i21_006,inst_doa_i21_005,inst_doa_i21_004,inst_doa_i21_003,inst_doa_i21_002,inst_doa_i21_001,inst_doa_i21_000}));
  // address_offset=22528;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'h0000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'h898989898A8A8A8A8A8A8B8B8B8B8B8B8C8C8C8C8C8C8D8D8D8D8D8D8D8E8E8E),
    .INIT_01(256'h8484848484858585858585858686868686868787878787878888888888888989),
    .INIT_02(256'h7F7F7F7F7F7F7F80808080808081818181818182828282828283838383838384),
    .INIT_03(256'h79797A7A7A7A7A7A7B7B7B7B7B7B7C7C7C7C7C7C7D7D7D7D7D7D7E7E7E7E7E7E),
    .INIT_04(256'h7474747575757575757676767676767777777777777878787878787979797979),
    .INIT_05(256'h6F6F6F6F70707070707071717171717172727272727273737373737374747474),
    .INIT_06(256'h6A6A6A6A6A6B6B6B6B6B6B6C6C6C6C6C6C6D6D6D6D6D6D6E6E6E6E6E6E6F6F6F),
    .INIT_07(256'h6565656565656666666666666767676767676868686868686969696969696A6A),
    .INIT_08(256'h6060606060606161616161616162626262626263636363636364646464646465),
    .INIT_09(256'h5A5B5B5B5B5B5B5C5C5C5C5C5C5D5D5D5D5D5D5D5E5E5E5E5E5E5F5F5F5F5F5F),
    .INIT_0A(256'h5555565656565656575757575757585858585858595959595959595A5A5A5A5A),
    .INIT_0B(256'h5050515151515151525252525252525353535353535454545454545555555555),
    .INIT_0C(256'h4B4B4B4C4C4C4C4C4C4D4D4D4D4D4D4E4E4E4E4E4E4E4F4F4F4F4F4F50505050),
    .INIT_0D(256'h464646474747474747484848484848484949494949494A4A4A4A4A4A4B4B4B4B),
    .INIT_0E(256'h4141414142424242424243434343434344444444444444454545454545464646),
    .INIT_0F(256'h3C3C3C3C3D3D3D3D3D3D3E3E3E3E3E3E3E3F3F3F3F3F3F404040404040414141),
    .INIT_10(256'h37373737383838383838383939393939393A3A3A3A3A3A3B3B3B3B3B3B3B3C3C),
    .INIT_11(256'h3232323233333333333333343434343434353535353535363636363636363737),
    .INIT_12(256'h2D2D2D2D2E2E2E2E2E2E2E2F2F2F2F2F2F303030303030303131313131313232),
    .INIT_13(256'h28282828282929292929292A2A2A2A2A2A2B2B2B2B2B2B2B2C2C2C2C2C2C2D2D),
    .INIT_14(256'h2323232324242424242424252525252525262626262626262727272727272828),
    .INIT_15(256'h1E1E1E1E1F1F1F1F1F1F1F202020202020212121212121212222222222222323),
    .INIT_16(256'h191919191A1A1A1A1A1A1A1B1B1B1B1B1B1C1C1C1C1C1C1C1D1D1D1D1D1D1E1E),
    .INIT_17(256'h1414141415151515151516161616161616171717171717181818181818181919),
    .INIT_18(256'h0F0F0F0F10101010101011111111111111121212121212131313131313141414),
    .INIT_19(256'h0A0A0A0B0B0B0B0B0B0B0C0C0C0C0C0C0D0D0D0D0D0D0D0E0E0E0E0E0E0F0F0F),
    .INIT_1A(256'h05050506060606060607070707070707080808080808090909090909090A0A0A),
    .INIT_1B(256'h0000010101010101010202020202020303030303030304040404040405050505),
    .INIT_1C(256'hFBFCFCFCFCFCFCFCFDFDFDFDFDFDFDFEFEFEFEFEFEFFFFFFFFFFFFFF00000000),
    .INIT_1D(256'hF6F7F7F7F7F7F7F8F8F8F8F8F8F8F9F9F9F9F9F9FAFAFAFAFAFAFAFBFBFBFBFB),
    .INIT_1E(256'hF2F2F2F2F2F2F3F3F3F3F3F3F3F4F4F4F4F4F4F4F5F5F5F5F5F5F6F6F6F6F6F6),
    .INIT_1F(256'hEDEDEDEDEDEDEEEEEEEEEEEEEFEFEFEFEFEFEFF0F0F0F0F0F0F1F1F1F1F1F1F1),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_022528_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_Naddra_o_al_n36 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i22_008,inst_doa_i22_007,inst_doa_i22_006,inst_doa_i22_005,inst_doa_i22_004,inst_doa_i22_003,inst_doa_i22_002,inst_doa_i22_001,inst_doa_i22_000}));
  // address_offset=23552;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hE8E8E8E8E8E9E9E9E9E9E9EAEAEAEAEAEAEAEBEBEBEBEBEBECECECECECECECED),
    .INIT_01(256'hE3E3E3E3E4E4E4E4E4E4E5E5E5E5E5E5E5E6E6E6E6E6E6E7E7E7E7E7E7E7E8E8),
    .INIT_02(256'hDEDEDFDFDFDFDFDFDFE0E0E0E0E0E0E0E1E1E1E1E1E1E2E2E2E2E2E2E2E3E3E3),
    .INIT_03(256'hD9DADADADADADADADBDBDBDBDBDBDCDCDCDCDCDCDCDDDDDDDDDDDDDDDEDEDEDE),
    .INIT_04(256'hD5D5D5D5D5D5D6D6D6D6D6D6D6D7D7D7D7D7D7D7D8D8D8D8D8D8D9D9D9D9D9D9),
    .INIT_05(256'hD0D0D0D0D0D1D1D1D1D1D1D1D2D2D2D2D2D2D3D3D3D3D3D3D3D4D4D4D4D4D4D4),
    .INIT_06(256'hCBCBCBCBCCCCCCCCCCCCCDCDCDCDCDCDCDCECECECECECECECFCFCFCFCFCFD0D0),
    .INIT_07(256'hC6C6C7C7C7C7C7C7C7C8C8C8C8C8C8C9C9C9C9C9C9C9CACACACACACACACBCBCB),
    .INIT_08(256'hC2C2C2C2C2C2C2C3C3C3C3C3C3C3C4C4C4C4C4C4C4C5C5C5C5C5C5C6C6C6C6C6),
    .INIT_09(256'hBDBDBDBDBDBEBEBEBEBEBEBEBFBFBFBFBFBFBFC0C0C0C0C0C0C0C1C1C1C1C1C1),
    .INIT_0A(256'hB8B8B8B9B9B9B9B9B9B9BABABABABABABABBBBBBBBBBBBBBBCBCBCBCBCBCBCBD),
    .INIT_0B(256'hB3B3B4B4B4B4B4B4B5B5B5B5B5B5B5B6B6B6B6B6B6B6B7B7B7B7B7B7B7B8B8B8),
    .INIT_0C(256'hAFAFAFAFAFAFB0B0B0B0B0B0B0B1B1B1B1B1B1B1B2B2B2B2B2B2B2B3B3B3B3B3),
    .INIT_0D(256'hAAAAAAAAABABABABABABABACACACACACACACADADADADADADADAEAEAEAEAEAEAF),
    .INIT_0E(256'hA5A5A6A6A6A6A6A6A6A7A7A7A7A7A7A7A8A8A8A8A8A8A9A9A9A9A9A9A9AAAAAA),
    .INIT_0F(256'hA1A1A1A1A1A1A2A2A2A2A2A2A2A3A3A3A3A3A3A3A4A4A4A4A4A4A4A5A5A5A5A5),
    .INIT_10(256'h9C9C9C9C9D9D9D9D9D9D9D9E9E9E9E9E9E9E9F9F9F9F9F9F9FA0A0A0A0A0A0A0),
    .INIT_11(256'h9797989898989898999999999999999A9A9A9A9A9A9A9B9B9B9B9B9B9B9C9C9C),
    .INIT_12(256'h9393939393939494949494949495959595959595969696969696969797979797),
    .INIT_13(256'h8E8E8E8F8F8F8F8F8F8F90909090909090919191919191919292929292929293),
    .INIT_14(256'h8A8A8A8A8A8A8A8B8B8B8B8B8B8B8C8C8C8C8C8C8C8D8D8D8D8D8D8D8E8E8E8E),
    .INIT_15(256'h8585858586868686868686878787878787878888888888888889898989898989),
    .INIT_16(256'h8081818181818181828282828282828383838383838384848484848484858585),
    .INIT_17(256'h7C7C7C7C7C7D7D7D7D7D7D7D7E7E7E7E7E7E7E7F7F7F7F7F7F7F808080808080),
    .INIT_18(256'h777778787878787878797979797979797A7A7A7A7A7A7A7B7B7B7B7B7B7B7C7C),
    .INIT_19(256'h7373737373737474747474747475757575757575767676767676767777777777),
    .INIT_1A(256'h6E6E6F6F6F6F6F6F6F6F70707070707070717171717171717272727272727273),
    .INIT_1B(256'h6A6A6A6A6A6A6B6B6B6B6B6B6B6C6C6C6C6C6C6C6D6D6D6D6D6D6D6E6E6E6E6E),
    .INIT_1C(256'h656566666666666666666767676767676768686868686868696969696969696A),
    .INIT_1D(256'h6161616161616262626262626263636363636363646464646464646565656565),
    .INIT_1E(256'h5C5C5D5D5D5D5D5D5D5E5E5E5E5E5E5E5F5F5F5F5F5F5F5F6060606060606061),
    .INIT_1F(256'h5858585858595959595959595A5A5A5A5A5A5A5A5B5B5B5B5B5B5B5C5C5C5C5C),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_023552_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_Naddra_o_al_n36 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i23_008,inst_doa_i23_007,inst_doa_i23_006,inst_doa_i23_005,inst_doa_i23_004,inst_doa_i23_003,inst_doa_i23_002,inst_doa_i23_001,inst_doa_i23_000}));
  // address_offset=24576;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'h5354545454545454555555555555555556565656565656575757575757575858),
    .INIT_01(256'h4F4F4F4F50505050505050505151515151515152525252525252535353535353),
    .INIT_02(256'h4B4B4B4B4B4B4B4C4C4C4C4C4C4C4C4D4D4D4D4D4D4D4E4E4E4E4E4E4E4F4F4F),
    .INIT_03(256'h464646474747474747474848484848484849494949494949494A4A4A4A4A4A4A),
    .INIT_04(256'h4242424242424343434343434344444444444444454545454545454546464646),
    .INIT_05(256'h3D3E3E3E3E3E3E3E3F3F3F3F3F3F3F3F40404040404040414141414141414242),
    .INIT_06(256'h393939393A3A3A3A3A3A3A3B3B3B3B3B3B3B3C3C3C3C3C3C3C3C3D3D3D3D3D3D),
    .INIT_07(256'h3535353535353636363636363637373737373737373838383838383839393939),
    .INIT_08(256'h3031313131313131313232323232323233333333333333343434343434343435),
    .INIT_09(256'h2C2C2C2D2D2D2D2D2D2D2D2E2E2E2E2E2E2E2F2F2F2F2F2F2F2F303030303030),
    .INIT_0A(256'h282828282828292929292929292A2A2A2A2A2A2A2A2B2B2B2B2B2B2B2C2C2C2C),
    .INIT_0B(256'h2424242424242424252525252525252626262626262626272727272727272828),
    .INIT_0C(256'h1F1F202020202020202021212121212121222222222222222223232323232323),
    .INIT_0D(256'h1B1B1B1B1C1C1C1C1C1C1C1C1D1D1D1D1D1D1D1E1E1E1E1E1E1E1E1F1F1F1F1F),
    .INIT_0E(256'h1717171717171818181818181818191919191919191A1A1A1A1A1A1A1A1B1B1B),
    .INIT_0F(256'h1313131313131313141414141414141515151515151515161616161616161617),
    .INIT_10(256'h0E0E0F0F0F0F0F0F0F1010101010101010111111111111111112121212121212),
    .INIT_11(256'h0A0A0A0B0B0B0B0B0B0B0B0C0C0C0C0C0C0C0C0D0D0D0D0D0D0D0E0E0E0E0E0E),
    .INIT_12(256'h060606060607070707070707080808080808080809090909090909090A0A0A0A),
    .INIT_13(256'h0202020202020303030303030303040404040404040505050505050505060606),
    .INIT_14(256'hFEFEFEFEFEFEFEFFFFFFFFFFFFFFFF0000000000000000010101010101010202),
    .INIT_15(256'hF9FAFAFAFAFAFAFAFBFBFBFBFBFBFBFBFCFCFCFCFCFCFCFCFDFDFDFDFDFDFDFD),
    .INIT_16(256'hF5F5F6F6F6F6F6F6F6F7F7F7F7F7F7F7F7F8F8F8F8F8F8F8F8F9F9F9F9F9F9F9),
    .INIT_17(256'hF1F1F1F2F2F2F2F2F2F2F3F3F3F3F3F3F3F3F4F4F4F4F4F4F4F4F5F5F5F5F5F5),
    .INIT_18(256'hEDEDEDEEEEEEEEEEEEEEEEEFEFEFEFEFEFEFEFF0F0F0F0F0F0F0F0F1F1F1F1F1),
    .INIT_19(256'hE9E9E9E9EAEAEAEAEAEAEAEAEBEBEBEBEBEBEBEBECECECECECECECEDEDEDEDED),
    .INIT_1A(256'hE5E5E5E5E6E6E6E6E6E6E6E6E7E7E7E7E7E7E7E7E8E8E8E8E8E8E8E8E9E9E9E9),
    .INIT_1B(256'hE1E1E1E1E1E2E2E2E2E2E2E2E2E3E3E3E3E3E3E3E3E4E4E4E4E4E4E4E4E5E5E5),
    .INIT_1C(256'hDDDDDDDDDDDEDEDEDEDEDEDEDEDFDFDFDFDFDFDFDFE0E0E0E0E0E0E0E0E1E1E1),
    .INIT_1D(256'hD9D9D9D9D9DADADADADADADADADBDBDBDBDBDBDBDBDCDCDCDCDCDCDCDCDDDDDD),
    .INIT_1E(256'hD5D5D5D5D5D6D6D6D6D6D6D6D6D7D7D7D7D7D7D7D7D8D8D8D8D8D8D8D8D9D9D9),
    .INIT_1F(256'hD1D1D1D1D1D2D2D2D2D2D2D2D2D3D3D3D3D3D3D3D3D4D4D4D4D4D4D4D4D5D5D5),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_024576_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_addra_o_al_n44 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i24_008,inst_doa_i24_007,inst_doa_i24_006,inst_doa_i24_005,inst_doa_i24_004,inst_doa_i24_003,inst_doa_i24_002,inst_doa_i24_001,inst_doa_i24_000}));
  // address_offset=24576;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'h0000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_024576_009 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n1580,open_n1581,open_n1582,open_n1583,open_n1584,open_n1585,open_n1586,1'b0,open_n1587}),
    .rsta(rsta),
    .doa({open_n1602,open_n1603,open_n1604,open_n1605,open_n1606,open_n1607,open_n1608,open_n1609,inst_doa_i24_009}));
  // address_offset=24576;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_024576_010 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n1638,open_n1639,open_n1640,open_n1641,open_n1642,open_n1643,open_n1644,1'b0,open_n1645}),
    .rsta(rsta),
    .doa({open_n1660,open_n1661,open_n1662,open_n1663,open_n1664,open_n1665,open_n1666,open_n1667,inst_doa_i24_010}));
  // address_offset=25600;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'hCDCDCDCDCDCECECECECECECECECFCFCFCFCFCFCFCFD0D0D0D0D0D0D0D0D1D1D1),
    .INIT_01(256'hC9C9C9C9C9CACACACACACACACACBCBCBCBCBCBCBCBCCCCCCCCCCCCCCCCCDCDCD),
    .INIT_02(256'hC5C5C5C5C5C6C6C6C6C6C6C6C6C7C7C7C7C7C7C7C7C8C8C8C8C8C8C8C8C9C9C9),
    .INIT_03(256'hC1C1C1C1C2C2C2C2C2C2C2C2C3C3C3C3C3C3C3C3C4C4C4C4C4C4C4C4C5C5C5C5),
    .INIT_04(256'hBDBDBDBEBEBEBEBEBEBEBEBEBFBFBFBFBFBFBFBFC0C0C0C0C0C0C0C0C1C1C1C1),
    .INIT_05(256'hB9B9B9BABABABABABABABABBBBBBBBBBBBBBBBBCBCBCBCBCBCBCBCBDBDBDBDBD),
    .INIT_06(256'hB5B5B6B6B6B6B6B6B6B6B7B7B7B7B7B7B7B7B8B8B8B8B8B8B8B8B9B9B9B9B9B9),
    .INIT_07(256'hB1B2B2B2B2B2B2B2B2B3B3B3B3B3B3B3B3B4B4B4B4B4B4B4B4B5B5B5B5B5B5B5),
    .INIT_08(256'hAEAEAEAEAEAEAEAEAFAFAFAFAFAFAFAFB0B0B0B0B0B0B0B0B1B1B1B1B1B1B1B1),
    .INIT_09(256'hAAAAAAAAAAAAABABABABABABABABABACACACACACACACACADADADADADADADADAE),
    .INIT_0A(256'hA6A6A6A6A6A7A7A7A7A7A7A7A7A8A8A8A8A8A8A8A8A8A9A9A9A9A9A9A9A9AAAA),
    .INIT_0B(256'hA2A2A2A2A3A3A3A3A3A3A3A3A4A4A4A4A4A4A4A4A5A5A5A5A5A5A5A5A5A6A6A6),
    .INIT_0C(256'h9E9E9F9F9F9F9F9F9F9FA0A0A0A0A0A0A0A0A0A1A1A1A1A1A1A1A1A2A2A2A2A2),
    .INIT_0D(256'h9B9B9B9B9B9B9B9B9C9C9C9C9C9C9C9C9C9D9D9D9D9D9D9D9D9E9E9E9E9E9E9E),
    .INIT_0E(256'h97979797979798989898989898989899999999999999999A9A9A9A9A9A9A9A9A),
    .INIT_0F(256'h9393939394949494949494949495959595959595959696969696969696969797),
    .INIT_10(256'h8F8F909090909090909090919191919191919192929292929292929293939393),
    .INIT_11(256'h8C8C8C8C8C8C8C8C8D8D8D8D8D8D8D8D8D8E8E8E8E8E8E8E8E8E8F8F8F8F8F8F),
    .INIT_12(256'h88888888888889898989898989898A8A8A8A8A8A8A8A8A8B8B8B8B8B8B8B8B8B),
    .INIT_13(256'h8484848585858585858585858686868686868686878787878787878787888888),
    .INIT_14(256'h8181818181818181818282828282828282828383838383838383848484848484),
    .INIT_15(256'h7D7D7D7D7D7D7E7E7E7E7E7E7E7E7E7F7F7F7F7F7F7F7F808080808080808080),
    .INIT_16(256'h7979797A7A7A7A7A7A7A7A7A7B7B7B7B7B7B7B7B7C7C7C7C7C7C7C7C7C7D7D7D),
    .INIT_17(256'h7676767676767676777777777777777777787878787878787878797979797979),
    .INIT_18(256'h7272727272737373737373737373747474747474747474757575757575757575),
    .INIT_19(256'h6E6F6F6F6F6F6F6F6F6F70707070707070707071717171717171717172727272),
    .INIT_1A(256'h6B6B6B6B6B6B6B6C6C6C6C6C6C6C6C6D6D6D6D6D6D6D6D6D6E6E6E6E6E6E6E6E),
    .INIT_1B(256'h6767676868686868686868686969696969696969696A6A6A6A6A6A6A6A6A6B6B),
    .INIT_1C(256'h6464646464646464656565656565656565666666666666666666676767676767),
    .INIT_1D(256'h6060606161616161616161616262626262626262626363636363636363636364),
    .INIT_1E(256'h5D5D5D5D5D5D5D5D5E5E5E5E5E5E5E5E5E5F5F5F5F5F5F5F5F5F606060606060),
    .INIT_1F(256'h5959595A5A5A5A5A5A5A5A5A5A5B5B5B5B5B5B5B5B5B5C5C5C5C5C5C5C5C5C5D),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_025600_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_addra_o_al_n44 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i25_008,inst_doa_i25_007,inst_doa_i25_006,inst_doa_i25_005,inst_doa_i25_004,inst_doa_i25_003,inst_doa_i25_002,inst_doa_i25_001,inst_doa_i25_000}));
  // address_offset=26624;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'h0000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'h5656565656565656575757575757575757585858585858585858595959595959),
    .INIT_01(256'h5252525353535353535353535454545454545454545455555555555555555556),
    .INIT_02(256'h4F4F4F4F4F4F4F50505050505050505050515151515151515151525252525252),
    .INIT_03(256'h4B4B4C4C4C4C4C4C4C4C4C4D4D4D4D4D4D4D4D4D4D4E4E4E4E4E4E4E4E4E4F4F),
    .INIT_04(256'h4848484848484949494949494949494A4A4A4A4A4A4A4A4A4A4B4B4B4B4B4B4B),
    .INIT_05(256'h4545454545454545454546464646464646464647474747474747474747484848),
    .INIT_06(256'h4141414142424242424242424243434343434343434343444444444444444444),
    .INIT_07(256'h3E3E3E3E3E3E3E3F3F3F3F3F3F3F3F3F3F404040404040404040414141414141),
    .INIT_08(256'h3A3B3B3B3B3B3B3B3B3B3B3C3C3C3C3C3C3C3C3C3D3D3D3D3D3D3D3D3D3D3E3E),
    .INIT_09(256'h3737373737383838383838383838393939393939393939393A3A3A3A3A3A3A3A),
    .INIT_0A(256'h3434343434343434353535353535353535363636363636363636363737373737),
    .INIT_0B(256'h3031313131313131313131323232323232323232333333333333333333333434),
    .INIT_0C(256'h2D2D2D2D2E2E2E2E2E2E2E2E2E2E2F2F2F2F2F2F2F2F2F303030303030303030),
    .INIT_0D(256'h2A2A2A2A2A2A2B2B2B2B2B2B2B2B2B2B2C2C2C2C2C2C2C2C2C2C2D2D2D2D2D2D),
    .INIT_0E(256'h27272727272727272728282828282828282828292929292929292929292A2A2A),
    .INIT_0F(256'h2324242424242424242424252525252525252525252626262626262626262627),
    .INIT_10(256'h2020202021212121212121212121222222222222222222222323232323232323),
    .INIT_11(256'h1D1D1D1D1D1D1E1E1E1E1E1E1E1E1E1E1F1F1F1F1F1F1F1F1F1F202020202020),
    .INIT_12(256'h1A1A1A1A1A1A1A1A1B1B1B1B1B1B1B1B1B1B1C1C1C1C1C1C1C1C1C1C1D1D1D1D),
    .INIT_13(256'h1717171717171717171818181818181818181818191919191919191919191A1A),
    .INIT_14(256'h1314141414141414141414151515151515151515151616161616161616161617),
    .INIT_15(256'h1010111111111111111111111112121212121212121212131313131313131313),
    .INIT_16(256'h0D0D0D0D0E0E0E0E0E0E0E0E0E0E0F0F0F0F0F0F0F0F0F0F1010101010101010),
    .INIT_17(256'h0A0A0A0A0A0B0B0B0B0B0B0B0B0B0B0C0C0C0C0C0C0C0C0C0C0D0D0D0D0D0D0D),
    .INIT_18(256'h07070707070708080808080808080808090909090909090909090A0A0A0A0A0A),
    .INIT_19(256'h0404040404040505050505050505050505060606060606060606060707070707),
    .INIT_1A(256'h0101010101010102020202020202020202020303030303030303030304040404),
    .INIT_1B(256'hFEFEFEFEFEFEFEFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000010101),
    .INIT_1C(256'hFBFBFBFBFBFBFBFBFCFCFCFCFCFCFCFCFCFCFDFDFDFDFDFDFDFDFDFDFDFEFEFE),
    .INIT_1D(256'hF8F8F8F8F8F8F8F8F9F9F9F9F9F9F9F9F9F9FAFAFAFAFAFAFAFAFAFAFAFBFBFB),
    .INIT_1E(256'hF5F5F5F5F5F5F5F5F6F6F6F6F6F6F6F6F6F6F7F7F7F7F7F7F7F7F7F7F7F8F8F8),
    .INIT_1F(256'hF2F2F2F2F2F2F2F3F3F3F3F3F3F3F3F3F3F3F4F4F4F4F4F4F4F4F4F4F4F5F5F5),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_026624_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_addra_o_al_n44 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i26_008,inst_doa_i26_007,inst_doa_i26_006,inst_doa_i26_005,inst_doa_i26_004,inst_doa_i26_003,inst_doa_i26_002,inst_doa_i26_001,inst_doa_i26_000}));
  // address_offset=27648;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hEFEFEFEFEFEFEFF0F0F0F0F0F0F0F0F0F0F0F1F1F1F1F1F1F1F1F1F1F1F2F2F2),
    .INIT_01(256'hECECECECECECEDEDEDEDEDEDEDEDEDEDEDEEEEEEEEEEEEEEEEEEEEEEEFEFEFEF),
    .INIT_02(256'hE9E9E9E9E9EAEAEAEAEAEAEAEAEAEAEAEBEBEBEBEBEBEBEBEBEBEBECECECECEC),
    .INIT_03(256'hE6E6E6E6E7E7E7E7E7E7E7E7E7E7E7E8E8E8E8E8E8E8E8E8E8E8E9E9E9E9E9E9),
    .INIT_04(256'hE3E3E3E4E4E4E4E4E4E4E4E4E4E4E5E5E5E5E5E5E5E5E5E5E5E6E6E6E6E6E6E6),
    .INIT_05(256'hE0E0E1E1E1E1E1E1E1E1E1E1E1E2E2E2E2E2E2E2E2E2E2E2E3E3E3E3E3E3E3E3),
    .INIT_06(256'hDEDEDEDEDEDEDEDEDEDEDEDFDFDFDFDFDFDFDFDFDFDFE0E0E0E0E0E0E0E0E0E0),
    .INIT_07(256'hDBDBDBDBDBDBDBDBDBDCDCDCDCDCDCDCDCDCDCDCDCDDDDDDDDDDDDDDDDDDDDDD),
    .INIT_08(256'hD8D8D8D8D8D8D8D9D9D9D9D9D9D9D9D9D9D9D9DADADADADADADADADADADADBDB),
    .INIT_09(256'hD5D5D5D5D5D6D6D6D6D6D6D6D6D6D6D6D6D7D7D7D7D7D7D7D7D7D7D7D8D8D8D8),
    .INIT_0A(256'hD2D2D2D3D3D3D3D3D3D3D3D3D3D3D4D4D4D4D4D4D4D4D4D4D4D4D5D5D5D5D5D5),
    .INIT_0B(256'hD0D0D0D0D0D0D0D0D0D0D0D0D1D1D1D1D1D1D1D1D1D1D1D2D2D2D2D2D2D2D2D2),
    .INIT_0C(256'hCDCDCDCDCDCDCDCDCDCECECECECECECECECECECECFCFCFCFCFCFCFCFCFCFCFCF),
    .INIT_0D(256'hCACACACACACACBCBCBCBCBCBCBCBCBCBCBCCCCCCCCCCCCCCCCCCCCCCCCCDCDCD),
    .INIT_0E(256'hC7C7C8C8C8C8C8C8C8C8C8C8C8C8C9C9C9C9C9C9C9C9C9C9C9C9CACACACACACA),
    .INIT_0F(256'hC5C5C5C5C5C5C5C5C5C5C6C6C6C6C6C6C6C6C6C6C6C6C7C7C7C7C7C7C7C7C7C7),
    .INIT_10(256'hC2C2C2C2C2C2C2C3C3C3C3C3C3C3C3C3C3C3C3C4C4C4C4C4C4C4C4C4C4C4C4C5),
    .INIT_11(256'hBFBFBFC0C0C0C0C0C0C0C0C0C0C0C0C1C1C1C1C1C1C1C1C1C1C1C1C2C2C2C2C2),
    .INIT_12(256'hBDBDBDBDBDBDBDBDBDBDBEBEBEBEBEBEBEBEBEBEBEBEBFBFBFBFBFBFBFBFBFBF),
    .INIT_13(256'hBABABABABABABBBBBBBBBBBBBBBBBBBBBBBBBCBCBCBCBCBCBCBCBCBCBCBCBDBD),
    .INIT_14(256'hB7B8B8B8B8B8B8B8B8B8B8B8B8B9B9B9B9B9B9B9B9B9B9B9B9B9BABABABABABA),
    .INIT_15(256'hB5B5B5B5B5B5B5B5B6B6B6B6B6B6B6B6B6B6B6B6B6B7B7B7B7B7B7B7B7B7B7B7),
    .INIT_16(256'hB2B2B2B3B3B3B3B3B3B3B3B3B3B3B3B3B4B4B4B4B4B4B4B4B4B4B4B4B5B5B5B5),
    .INIT_17(256'hB0B0B0B0B0B0B0B0B0B0B1B1B1B1B1B1B1B1B1B1B1B1B1B2B2B2B2B2B2B2B2B2),
    .INIT_18(256'hADADADADAEAEAEAEAEAEAEAEAEAEAEAEAEAFAFAFAFAFAFAFAFAFAFAFAFAFB0B0),
    .INIT_19(256'hABABABABABABABABABABABACACACACACACACACACACACACACADADADADADADADAD),
    .INIT_1A(256'hA8A8A8A8A8A9A9A9A9A9A9A9A9A9A9A9A9AAAAAAAAAAAAAAAAAAAAAAAAAAABAB),
    .INIT_1B(256'hA6A6A6A6A6A6A6A6A6A6A6A7A7A7A7A7A7A7A7A7A7A7A7A7A8A8A8A8A8A8A8A8),
    .INIT_1C(256'hA3A3A3A3A4A4A4A4A4A4A4A4A4A4A4A4A4A5A5A5A5A5A5A5A5A5A5A5A5A5A6A6),
    .INIT_1D(256'hA1A1A1A1A1A1A1A1A1A1A2A2A2A2A2A2A2A2A2A2A2A2A2A3A3A3A3A3A3A3A3A3),
    .INIT_1E(256'h9E9E9E9F9F9F9F9F9F9F9F9F9F9F9F9FA0A0A0A0A0A0A0A0A0A0A0A0A0A1A1A1),
    .INIT_1F(256'h9C9C9C9C9C9C9C9C9D9D9D9D9D9D9D9D9D9D9D9D9D9E9E9E9E9E9E9E9E9E9E9E),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_027648_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_addra_o_al_n44 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i27_008,inst_doa_i27_007,inst_doa_i27_006,inst_doa_i27_005,inst_doa_i27_004,inst_doa_i27_003,inst_doa_i27_002,inst_doa_i27_001,inst_doa_i27_000}));
  // address_offset=28672;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h9A9A9A9A9A9A9A9A9A9A9A9A9A9B9B9B9B9B9B9B9B9B9B9B9B9B9B9C9C9C9C9C),
    .INIT_01(256'h9797979797989898989898989898989898989899999999999999999999999999),
    .INIT_02(256'h9595959595959595959596969696969696969696969696969797979797979797),
    .INIT_03(256'h9293939393939393939393939393939494949494949494949494949495959595),
    .INIT_04(256'h9090909090909191919191919191919191919192929292929292929292929292),
    .INIT_05(256'h8E8E8E8E8E8E8E8E8E8E8F8F8F8F8F8F8F8F8F8F8F8F8F8F9090909090909090),
    .INIT_06(256'h8C8C8C8C8C8C8C8C8C8C8C8C8C8C8D8D8D8D8D8D8D8D8D8D8D8D8D8D8E8E8E8E),
    .INIT_07(256'h898989898A8A8A8A8A8A8A8A8A8A8A8A8A8A8B8B8B8B8B8B8B8B8B8B8B8B8B8B),
    .INIT_08(256'h8787878787878788888888888888888888888888888889898989898989898989),
    .INIT_09(256'h8585858585858585858585868686868686868686868686868687878787878787),
    .INIT_0A(256'h8383838383838383838383838383848484848484848484848484848485858585),
    .INIT_0B(256'h8080818181818181818181818181818181828282828282828282828282828282),
    .INIT_0C(256'h7E7E7E7E7E7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F808080808080808080808080),
    .INIT_0D(256'h7C7C7C7C7C7C7C7C7D7D7D7D7D7D7D7D7D7D7D7D7D7D7E7E7E7E7E7E7E7E7E7E),
    .INIT_0E(256'h7A7A7A7A7A7A7A7A7A7A7B7B7B7B7B7B7B7B7B7B7B7B7B7B7B7C7C7C7C7C7C7C),
    .INIT_0F(256'h7878787878787878787878787979797979797979797979797979797A7A7A7A7A),
    .INIT_10(256'h7676767676767676767676767677777777777777777777777777777777787878),
    .INIT_11(256'h7474747474747474747474747474747575757575757575757575757575757676),
    .INIT_12(256'h7172727272727272727272727272727273737373737373737373737373737373),
    .INIT_13(256'h6F6F707070707070707070707070707070717171717171717171717171717171),
    .INIT_14(256'h6D6D6E6E6E6E6E6E6E6E6E6E6E6E6E6E6E6E6F6F6F6F6F6F6F6F6F6F6F6F6F6F),
    .INIT_15(256'h6B6B6C6C6C6C6C6C6C6C6C6C6C6C6C6C6C6C6D6D6D6D6D6D6D6D6D6D6D6D6D6D),
    .INIT_16(256'h69696A6A6A6A6A6A6A6A6A6A6A6A6A6A6A6A6B6B6B6B6B6B6B6B6B6B6B6B6B6B),
    .INIT_17(256'h6767686868686868686868686868686868686969696969696969696969696969),
    .INIT_18(256'h6566666666666666666666666666666666666767676767676767676767676767),
    .INIT_19(256'h6364646464646464646464646464646464656565656565656565656565656565),
    .INIT_1A(256'h6262626262626262626262626262626263636363636363636363636363636363),
    .INIT_1B(256'h6060606060606060606060606060606161616161616161616161616161616162),
    .INIT_1C(256'h5E5E5E5E5E5E5E5E5E5E5E5E5E5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F6060),
    .INIT_1D(256'h5C5C5C5C5C5C5C5C5C5C5C5D5D5D5D5D5D5D5D5D5D5D5D5D5D5D5D5D5E5E5E5E),
    .INIT_1E(256'h5A5A5A5A5A5A5A5A5B5B5B5B5B5B5B5B5B5B5B5B5B5B5B5B5B5B5C5C5C5C5C5C),
    .INIT_1F(256'h58585858585959595959595959595959595959595959595A5A5A5A5A5A5A5A5A),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_028672_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_addra[_o_al_n52 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i28_008,inst_doa_i28_007,inst_doa_i28_006,inst_doa_i28_005,inst_doa_i28_004,inst_doa_i28_003,inst_doa_i28_002,inst_doa_i28_001,inst_doa_i28_000}));
  // address_offset=29696;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h5656575757575757575757575757575757575757585858585858585858585858),
    .INIT_01(256'h5555555555555555555555555555555556565656565656565656565656565656),
    .INIT_02(256'h5353535353535353535353535354545454545454545454545454545454545455),
    .INIT_03(256'h5151515151515151525252525252525252525252525252525252535353535353),
    .INIT_04(256'h4F4F4F4F50505050505050505050505050505050505051515151515151515151),
    .INIT_05(256'h4E4E4E4E4E4E4E4E4E4E4E4E4E4E4E4E4E4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F),
    .INIT_06(256'h4C4C4C4C4C4C4C4C4C4C4C4C4D4D4D4D4D4D4D4D4D4D4D4D4D4D4D4D4D4D4E4E),
    .INIT_07(256'h4A4A4A4A4A4A4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4C4C4C4C4C4C4C),
    .INIT_08(256'h494949494949494949494949494949494949494A4A4A4A4A4A4A4A4A4A4A4A4A),
    .INIT_09(256'h4747474747474747474747474848484848484848484848484848484848484849),
    .INIT_0A(256'h4545454545464646464646464646464646464646464646464647474747474747),
    .INIT_0B(256'h4444444444444444444444444444444444454545454545454545454545454545),
    .INIT_0C(256'h4242424242424242424343434343434343434343434343434343434343444444),
    .INIT_0D(256'h4041414141414141414141414141414141414141414242424242424242424242),
    .INIT_0E(256'h3F3F3F3F3F3F3F3F3F3F3F3F4040404040404040404040404040404040404040),
    .INIT_0F(256'h3D3D3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3F3F3F3F3F3F3F3F3F),
    .INIT_10(256'h3C3C3C3C3C3C3C3C3C3C3C3C3C3D3D3D3D3D3D3D3D3D3D3D3D3D3D3D3D3D3D3D),
    .INIT_11(256'h3A3A3A3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3C3C3C3C3C3C3C3C),
    .INIT_12(256'h393939393939393939393939393A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A),
    .INIT_13(256'h3737383838383838383838383838383838383838383838383939393939393939),
    .INIT_14(256'h3636363636363636363636373737373737373737373737373737373737373737),
    .INIT_15(256'h3535353535353535353535353535353535353535353636363636363636363636),
    .INIT_16(256'h3333333333333333343434343434343434343434343434343434343434343435),
    .INIT_17(256'h3232323232323232323232323232323232333333333333333333333333333333),
    .INIT_18(256'h3030313131313131313131313131313131313131313131313131323232323232),
    .INIT_19(256'h2F2F2F2F2F2F2F2F2F2F2F303030303030303030303030303030303030303030),
    .INIT_1A(256'h2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2F2F2F2F2F2F2F2F2F2F2F2F2F),
    .INIT_1B(256'h2C2C2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2E2E2E2E2E),
    .INIT_1C(256'h2B2B2B2B2B2B2B2B2B2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C),
    .INIT_1D(256'h2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B),
    .INIT_1E(256'h29292929292929292929292929292929292929292929292A2A2A2A2A2A2A2A2A),
    .INIT_1F(256'h2727272728282828282828282828282828282828282828282828282828282929),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_029696_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_addra[_o_al_n52 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i29_008,inst_doa_i29_007,inst_doa_i29_006,inst_doa_i29_005,inst_doa_i29_004,inst_doa_i29_003,inst_doa_i29_002,inst_doa_i29_001,inst_doa_i29_000}));
  // address_offset=30720;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h2626262626262626262727272727272727272727272727272727272727272727),
    .INIT_01(256'h2525252525252525252525252525252626262626262626262626262626262626),
    .INIT_02(256'h2424242424242424242424242424242424242424252525252525252525252525),
    .INIT_03(256'h2323232323232323232323232323232323232323232323232324242424242424),
    .INIT_04(256'h2122222222222222222222222222222222222222222222222222222222232323),
    .INIT_05(256'h2020202021212121212121212121212121212121212121212121212121212121),
    .INIT_06(256'h1F1F1F1F1F1F1F20202020202020202020202020202020202020202020202020),
    .INIT_07(256'h1E1E1E1E1E1E1E1E1E1E1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F),
    .INIT_08(256'h1D1D1D1D1D1D1D1D1D1D1D1D1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E),
    .INIT_09(256'h1C1C1C1C1C1C1C1C1C1C1C1C1C1C1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D),
    .INIT_0A(256'h1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C),
    .INIT_0B(256'h1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B),
    .INIT_0C(256'h1919191919191919191919191919191A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A),
    .INIT_0D(256'h1818181818181818181818181818181919191919191919191919191919191919),
    .INIT_0E(256'h1717171717171717171717171718181818181818181818181818181818181818),
    .INIT_0F(256'h1616161616161616161616171717171717171717171717171717171717171717),
    .INIT_10(256'h1515151515151515161616161616161616161616161616161616161616161616),
    .INIT_11(256'h1414141414151515151515151515151515151515151515151515151515151515),
    .INIT_12(256'h1414141414141414141414141414141414141414141414141414141414141414),
    .INIT_13(256'h1313131313131313131313131313131313131313131313131313131313131313),
    .INIT_14(256'h1212121212121212121212121212121212121212121212121212121313131313),
    .INIT_15(256'h1111111111111111111111111111111111111111121212121212121212121212),
    .INIT_16(256'h1010101010101010101010101011111111111111111111111111111111111111),
    .INIT_17(256'h0F0F0F0F10101010101010101010101010101010101010101010101010101010),
    .INIT_18(256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F),
    .INIT_19(256'h0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0F0F0F0F0F0F),
    .INIT_1A(256'h0D0D0D0D0D0D0D0D0D0D0D0D0D0D0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E),
    .INIT_1B(256'h0C0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D),
    .INIT_1C(256'h0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C),
    .INIT_1D(256'h0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0C0C0C0C0C0C0C0C0C0C0C0C0C0C),
    .INIT_1E(256'h0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B),
    .INIT_1F(256'h0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_030720_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_addra[_o_al_n52 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i30_008,inst_doa_i30_007,inst_doa_i30_006,inst_doa_i30_005,inst_doa_i30_004,inst_doa_i30_003,inst_doa_i30_002,inst_doa_i30_001,inst_doa_i30_000}));
  // address_offset=31744;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h090909090909090909090909090A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A),
    .INIT_01(256'h0909090909090909090909090909090909090909090909090909090909090909),
    .INIT_02(256'h0808080808080808080808080808080808080808080809090909090909090909),
    .INIT_03(256'h0808080808080808080808080808080808080808080808080808080808080808),
    .INIT_04(256'h0707070707070707070707070707070707070707070707070707070707080808),
    .INIT_05(256'h0707070707070707070707070707070707070707070707070707070707070707),
    .INIT_06(256'h0606060606060606060606060606060606060606060606060606060606060607),
    .INIT_07(256'h0606060606060606060606060606060606060606060606060606060606060606),
    .INIT_08(256'h0505050505050505050505050505050505050505050505050505050506060606),
    .INIT_09(256'h0505050505050505050505050505050505050505050505050505050505050505),
    .INIT_0A(256'h0404040404040404040404040404040404040405050505050505050505050505),
    .INIT_0B(256'h0404040404040404040404040404040404040404040404040404040404040404),
    .INIT_0C(256'h0304040404040404040404040404040404040404040404040404040404040404),
    .INIT_0D(256'h0303030303030303030303030303030303030303030303030303030303030303),
    .INIT_0E(256'h0303030303030303030303030303030303030303030303030303030303030303),
    .INIT_0F(256'h0202020303030303030303030303030303030303030303030303030303030303),
    .INIT_10(256'h0202020202020202020202020202020202020202020202020202020202020202),
    .INIT_11(256'h0202020202020202020202020202020202020202020202020202020202020202),
    .INIT_12(256'h0202020202020202020202020202020202020202020202020202020202020202),
    .INIT_13(256'h0101010101010101010101010101010202020202020202020202020202020202),
    .INIT_14(256'h0101010101010101010101010101010101010101010101010101010101010101),
    .INIT_15(256'h0101010101010101010101010101010101010101010101010101010101010101),
    .INIT_16(256'h0101010101010101010101010101010101010101010101010101010101010101),
    .INIT_17(256'h0101010101010101010101010101010101010101010101010101010101010101),
    .INIT_18(256'h0000000000000101010101010101010101010101010101010101010101010101),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_031744_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_addra[_o_al_n52 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i31_008,inst_doa_i31_007,inst_doa_i31_006,inst_doa_i31_005,inst_doa_i31_004,inst_doa_i31_003,inst_doa_i31_002,inst_doa_i31_001,inst_doa_i31_000}));
  // address_offset=32768;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0101010101010101010101010101010101010101010101010100000000000000),
    .INIT_08(256'h0101010101010101010101010101010101010101010101010101010101010101),
    .INIT_09(256'h0101010101010101010101010101010101010101010101010101010101010101),
    .INIT_0A(256'h0101010101010101010101010101010101010101010101010101010101010101),
    .INIT_0B(256'h0101010101010101010101010101010101010101010101010101010101010101),
    .INIT_0C(256'h0202020202020202020202020202020201010101010101010101010101010101),
    .INIT_0D(256'h0202020202020202020202020202020202020202020202020202020202020202),
    .INIT_0E(256'h0202020202020202020202020202020202020202020202020202020202020202),
    .INIT_0F(256'h0202020202020202020202020202020202020202020202020202020202020202),
    .INIT_10(256'h0303030303030303030303030303030303030303030303030303030302020202),
    .INIT_11(256'h0303030303030303030303030303030303030303030303030303030303030303),
    .INIT_12(256'h0303030303030303030303030303030303030303030303030303030303030303),
    .INIT_13(256'h0404040404040404040404040404040404040404040404040404040404040303),
    .INIT_14(256'h0404040404040404040404040404040404040404040404040404040404040404),
    .INIT_15(256'h0505050505050505050505050404040404040404040404040404040404040404),
    .INIT_16(256'h0505050505050505050505050505050505050505050505050505050505050505),
    .INIT_17(256'h0606060505050505050505050505050505050505050505050505050505050505),
    .INIT_18(256'h0606060606060606060606060606060606060606060606060606060606060606),
    .INIT_19(256'h0606060606060606060606060606060606060606060606060606060606060606),
    .INIT_1A(256'h0707070707070707070707070707070707070707070707070707070707070707),
    .INIT_1B(256'h0808070707070707070707070707070707070707070707070707070707070707),
    .INIT_1C(256'h0808080808080808080808080808080808080808080808080808080808080808),
    .INIT_1D(256'h0909090909090909090808080808080808080808080808080808080808080808),
    .INIT_1E(256'h0909090909090909090909090909090909090909090909090909090909090909),
    .INIT_1F(256'h0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0909090909090909090909090909),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_032768_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_Naddr_o_al_n60 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i32_008,inst_doa_i32_007,inst_doa_i32_006,inst_doa_i32_005,inst_doa_i32_004,inst_doa_i32_003,inst_doa_i32_002,inst_doa_i32_001,inst_doa_i32_000}));
  // address_offset=32768;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000000000000000),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_032768_009 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n2032,open_n2033,open_n2034,open_n2035,open_n2036,open_n2037,open_n2038,1'b0,open_n2039}),
    .rsta(rsta),
    .doa({open_n2054,open_n2055,open_n2056,open_n2057,open_n2058,open_n2059,open_n2060,open_n2061,inst_doa_i32_009}));
  // address_offset=32768;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_032768_010 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n2090,open_n2091,open_n2092,open_n2093,open_n2094,open_n2095,open_n2096,1'b0,open_n2097}),
    .rsta(rsta),
    .doa({open_n2112,open_n2113,open_n2114,open_n2115,open_n2116,open_n2117,open_n2118,open_n2119,inst_doa_i32_010}));
  // address_offset=33792;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A),
    .INIT_01(256'h0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0A),
    .INIT_02(256'h0C0C0C0C0C0C0C0C0C0C0C0C0C0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0B),
    .INIT_03(256'h0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C),
    .INIT_04(256'h0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D0C0C),
    .INIT_05(256'h0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0D0D0D0D0D0D0D0D0D0D0D0D0D0D0D),
    .INIT_06(256'h0F0F0F0F0F0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E),
    .INIT_07(256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F),
    .INIT_08(256'h1010101010101010101010101010101010101010101010101010100F0F0F0F0F),
    .INIT_09(256'h1111111111111111111111111111111111111010101010101010101010101010),
    .INIT_0A(256'h1212121212121212121212111111111111111111111111111111111111111111),
    .INIT_0B(256'h1313131312121212121212121212121212121212121212121212121212121212),
    .INIT_0C(256'h1313131313131313131313131313131313131313131313131313131313131313),
    .INIT_0D(256'h1414141414141414141414141414141414141414141414141414141414141413),
    .INIT_0E(256'h1515151515151515151515151515151515151515151515151515141414141414),
    .INIT_0F(256'h1616161616161616161616161616161616161616161616151515151515151515),
    .INIT_10(256'h1717171717171717171717171717171717171717161616161616161616161616),
    .INIT_11(256'h1818181818181818181818181818181818181717171717171717171717171717),
    .INIT_12(256'h1919191919191919191919191919191918181818181818181818181818181818),
    .INIT_13(256'h1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A19191919191919191919191919191919),
    .INIT_14(256'h1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A1A),
    .INIT_15(256'h1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B),
    .INIT_16(256'h1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C),
    .INIT_17(256'h1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1D1D1D1D1D1D1D1D1D1D1D1D1D),
    .INIT_18(256'h1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1E1E1E1E1E1E1E1E1E1E1E),
    .INIT_19(256'h2020202020202020202020202020202020202020202020201F1F1F1F1F1F1F1F),
    .INIT_1A(256'h2121212121212121212121212121212121212121212121212121212020202020),
    .INIT_1B(256'h2323222222222222222222222222222222222222222222222222222222222121),
    .INIT_1C(256'h2424242424242323232323232323232323232323232323232323232323232323),
    .INIT_1D(256'h2525252525252525252525242424242424242424242424242424242424242424),
    .INIT_1E(256'h2626262626262626262626262626262625252525252525252525252525252525),
    .INIT_1F(256'h2727272727272727272727272727272727272727272726262626262626262626),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_033792_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_Naddr_o_al_n60 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i33_008,inst_doa_i33_007,inst_doa_i33_006,inst_doa_i33_005,inst_doa_i33_004,inst_doa_i33_003,inst_doa_i33_002,inst_doa_i33_001,inst_doa_i33_000}));
  // address_offset=34816;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h2928282828282828282828282828282828282828282828282828282727272727),
    .INIT_01(256'h2A2A2A2A2A2A2A2A292929292929292929292929292929292929292929292929),
    .INIT_02(256'h2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A),
    .INIT_03(256'h2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2B2B2B2B2B2B2B2B2B2B),
    .INIT_04(256'h2E2E2E2E2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2C2C2C),
    .INIT_05(256'h2F2F2F2F2F2F2F2F2F2F2F2F2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E),
    .INIT_06(256'h30303030303030303030303030303030303030302F2F2F2F2F2F2F2F2F2F2F2F),
    .INIT_07(256'h3232323232313131313131313131313131313131313131313131313131303030),
    .INIT_08(256'h3333333333333333333333333333323232323232323232323232323232323232),
    .INIT_09(256'h3434343434343434343434343434343434343434343434333333333333333333),
    .INIT_0A(256'h3636363636363636363635353535353535353535353535353535353535353535),
    .INIT_0B(256'h3737373737373737373737373737373737373737363636363636363636363636),
    .INIT_0C(256'h3939393939393938383838383838383838383838383838383838383838373737),
    .INIT_0D(256'h3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3A3939393939393939393939393939),
    .INIT_0E(256'h3C3C3C3C3C3C3C3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3B3A3A3A3A),
    .INIT_0F(256'h3D3D3D3D3D3D3D3D3D3D3D3D3D3D3D3D3D3D3C3C3C3C3C3C3C3C3C3C3C3C3C3C),
    .INIT_10(256'h3F3F3F3F3F3F3F3F3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3D3D3D),
    .INIT_11(256'h404040404040404040404040404040404040403F3F3F3F3F3F3F3F3F3F3F3F3F),
    .INIT_12(256'h4242424242424242424241414141414141414141414141414141414141414040),
    .INIT_13(256'h4444434343434343434343434343434343434343434342424242424242424242),
    .INIT_14(256'h4545454545454545454545454545444444444444444444444444444444444444),
    .INIT_15(256'h4747474747474646464646464646464646464646464646464646454545454545),
    .INIT_16(256'h4848484848484848484848484848484848484847474747474747474747474747),
    .INIT_17(256'h4A4A4A4A4A4A4A4A4A4A4A4A4949494949494949494949494949494949494949),
    .INIT_18(256'h4C4C4C4C4C4C4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4A4A4A4A4A4A4A),
    .INIT_19(256'h4E4D4D4D4D4D4D4D4D4D4D4D4D4D4D4D4D4D4D4C4C4C4C4C4C4C4C4C4C4C4C4C),
    .INIT_1A(256'h4F4F4F4F4F4F4F4F4F4F4F4F4F4F4E4E4E4E4E4E4E4E4E4E4E4E4E4E4E4E4E4E),
    .INIT_1B(256'h5151515151515151515050505050505050505050505050505050504F4F4F4F4F),
    .INIT_1C(256'h5353535353525252525252525252525252525252525252515151515151515151),
    .INIT_1D(256'h5454545454545454545454545454545454545353535353535353535353535353),
    .INIT_1E(256'h5656565656565656565656565656565555555555555555555555555555555555),
    .INIT_1F(256'h5858585858585858585858575757575757575757575757575757575757565656),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_034816_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_Naddr_o_al_n60 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i34_008,inst_doa_i34_007,inst_doa_i34_006,inst_doa_i34_005,inst_doa_i34_004,inst_doa_i34_003,inst_doa_i34_002,inst_doa_i34_001,inst_doa_i34_000}));
  // address_offset=35840;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h5A5A5A5A5A5A5A5A595959595959595959595959595959595959585858585858),
    .INIT_01(256'h5C5C5C5C5C5C5B5B5B5B5B5B5B5B5B5B5B5B5B5B5B5B5B5A5A5A5A5A5A5A5A5A),
    .INIT_02(256'h5E5E5E5D5D5D5D5D5D5D5D5D5D5D5D5D5D5D5D5D5C5C5C5C5C5C5C5C5C5C5C5C),
    .INIT_03(256'h605F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5E5E5E5E5E5E5E5E5E5E5E5E5E5E),
    .INIT_04(256'h6161616161616161616161616161616160606060606060606060606060606060),
    .INIT_05(256'h6363636363636363636363636363636262626262626262626262626262626262),
    .INIT_06(256'h6565656565656565656565656565646464646464646464646464646464646363),
    .INIT_07(256'h6767676767676767676767676766666666666666666666666666666666666565),
    .INIT_08(256'h6969696969696969696969696968686868686868686868686868686868676767),
    .INIT_09(256'h6B6B6B6B6B6B6B6B6B6B6B6B6B6A6A6A6A6A6A6A6A6A6A6A6A6A6A6A6A696969),
    .INIT_0A(256'h6D6D6D6D6D6D6D6D6D6D6D6D6D6C6C6C6C6C6C6C6C6C6C6C6C6C6C6C6C6B6B6B),
    .INIT_0B(256'h6F6F6F6F6F6F6F6F6F6F6F6F6F6E6E6E6E6E6E6E6E6E6E6E6E6E6E6E6E6D6D6D),
    .INIT_0C(256'h71717171717171717171717171717070707070707070707070707070706F6F6F),
    .INIT_0D(256'h7373737373737373737373737373737272727272727272727272727272727171),
    .INIT_0E(256'h7675757575757575757575757575757574747474747474747474747474747473),
    .INIT_0F(256'h7878777777777777777777777777777777777676767676767676767676767676),
    .INIT_10(256'h7A7A7A7A79797979797979797979797979797978787878787878787878787878),
    .INIT_11(256'h7C7C7C7C7C7C7B7B7B7B7B7B7B7B7B7B7B7B7B7B7B7A7A7A7A7A7A7A7A7A7A7A),
    .INIT_12(256'h7E7E7E7E7E7E7E7E7E7D7D7D7D7D7D7D7D7D7D7D7D7D7D7C7C7C7C7C7C7C7C7C),
    .INIT_13(256'h80808080808080808080807F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7E7E7E7E7E7E),
    .INIT_14(256'h8282828282828282828282828282818181818181818181818181818181808080),
    .INIT_15(256'h8585858484848484848484848484848484838383838383838383838383838382),
    .INIT_16(256'h8787878787878686868686868686868686868686858585858585858585858585),
    .INIT_17(256'h8989898989898989898888888888888888888888888888888787878787878787),
    .INIT_18(256'h8B8B8B8B8B8B8B8B8B8B8B8B8B8A8A8A8A8A8A8A8A8A8A8A8A8A8A8989898989),
    .INIT_19(256'h8E8E8E8D8D8D8D8D8D8D8D8D8D8D8D8D8D8C8C8C8C8C8C8C8C8C8C8C8C8C8C8B),
    .INIT_1A(256'h909090909090908F8F8F8F8F8F8F8F8F8F8F8F8F8F8E8E8E8E8E8E8E8E8E8E8E),
    .INIT_1B(256'h9292929292929292929292929191919191919191919191919190909090909090),
    .INIT_1C(256'h9595959494949494949494949494949493939393939393939393939393939292),
    .INIT_1D(256'h9797979797979796969696969696969696969696969595959595959595959595),
    .INIT_1E(256'h9999999999999999999999999898989898989898989898989898979797979797),
    .INIT_1F(256'h9C9C9C9C9B9B9B9B9B9B9B9B9B9B9B9B9B9B9A9A9A9A9A9A9A9A9A9A9A9A9A99),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_035840_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_Naddr_o_al_n60 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i35_008,inst_doa_i35_007,inst_doa_i35_006,inst_doa_i35_005,inst_doa_i35_004,inst_doa_i35_003,inst_doa_i35_002,inst_doa_i35_001,inst_doa_i35_000}));
  // address_offset=36864;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h9E9E9E9E9E9E9E9E9E9E9D9D9D9D9D9D9D9D9D9D9D9D9D9C9C9C9C9C9C9C9C9C),
    .INIT_01(256'hA1A1A0A0A0A0A0A0A0A0A0A0A0A0A09F9F9F9F9F9F9F9F9F9F9F9F9F9E9E9E9E),
    .INIT_02(256'hA3A3A3A3A3A3A3A3A2A2A2A2A2A2A2A2A2A2A2A2A2A1A1A1A1A1A1A1A1A1A1A1),
    .INIT_03(256'hA6A5A5A5A5A5A5A5A5A5A5A5A5A5A4A4A4A4A4A4A4A4A4A4A4A4A4A3A3A3A3A3),
    .INIT_04(256'hA8A8A8A8A8A8A8A7A7A7A7A7A7A7A7A7A7A7A7A7A6A6A6A6A6A6A6A6A6A6A6A6),
    .INIT_05(256'hABAAAAAAAAAAAAAAAAAAAAAAAAAAA9A9A9A9A9A9A9A9A9A9A9A9A8A8A8A8A8A8),
    .INIT_06(256'hADADADADADADADACACACACACACACACACACACACACABABABABABABABABABABABAB),
    .INIT_07(256'hB0AFAFAFAFAFAFAFAFAFAFAFAFAFAEAEAEAEAEAEAEAEAEAEAEAEAEADADADADAD),
    .INIT_08(256'hB2B2B2B2B2B2B2B2B1B1B1B1B1B1B1B1B1B1B1B1B1B0B0B0B0B0B0B0B0B0B0B0),
    .INIT_09(256'hB5B5B5B4B4B4B4B4B4B4B4B4B4B4B4B3B3B3B3B3B3B3B3B3B3B3B3B3B2B2B2B2),
    .INIT_0A(256'hB7B7B7B7B7B7B7B7B7B7B6B6B6B6B6B6B6B6B6B6B6B6B6B5B5B5B5B5B5B5B5B5),
    .INIT_0B(256'hBABABABABAB9B9B9B9B9B9B9B9B9B9B9B9B9B8B8B8B8B8B8B8B8B8B8B8B8B7B7),
    .INIT_0C(256'hBDBCBCBCBCBCBCBCBCBCBCBCBCBBBBBBBBBBBBBBBBBBBBBBBBBABABABABABABA),
    .INIT_0D(256'hBFBFBFBFBFBFBFBFBFBEBEBEBEBEBEBEBEBEBEBEBEBDBDBDBDBDBDBDBDBDBDBD),
    .INIT_0E(256'hC2C2C2C2C1C1C1C1C1C1C1C1C1C1C1C1C0C0C0C0C0C0C0C0C0C0C0C0BFBFBFBF),
    .INIT_0F(256'hC4C4C4C4C4C4C4C4C4C4C4C4C3C3C3C3C3C3C3C3C3C3C3C3C2C2C2C2C2C2C2C2),
    .INIT_10(256'hC7C7C7C7C7C7C7C7C7C6C6C6C6C6C6C6C6C6C6C6C6C5C5C5C5C5C5C5C5C5C5C5),
    .INIT_11(256'hCACACACACAC9C9C9C9C9C9C9C9C9C9C9C9C8C8C8C8C8C8C8C8C8C8C8C8C7C7C7),
    .INIT_12(256'hCDCDCCCCCCCCCCCCCCCCCCCCCCCCCBCBCBCBCBCBCBCBCBCBCBCACACACACACACA),
    .INIT_13(256'hCFCFCFCFCFCFCFCFCFCFCFCECECECECECECECECECECECDCDCDCDCDCDCDCDCDCD),
    .INIT_14(256'hD2D2D2D2D2D2D2D2D1D1D1D1D1D1D1D1D1D1D1D0D0D0D0D0D0D0D0D0D0D0D0CF),
    .INIT_15(256'hD5D5D5D5D5D4D4D4D4D4D4D4D4D4D4D4D4D3D3D3D3D3D3D3D3D3D3D3D2D2D2D2),
    .INIT_16(256'hD8D8D8D7D7D7D7D7D7D7D7D7D7D7D6D6D6D6D6D6D6D6D6D6D6D6D5D5D5D5D5D5),
    .INIT_17(256'hDBDADADADADADADADADADADAD9D9D9D9D9D9D9D9D9D9D9D9D8D8D8D8D8D8D8D8),
    .INIT_18(256'hDDDDDDDDDDDDDDDDDDDDDCDCDCDCDCDCDCDCDCDCDCDCDBDBDBDBDBDBDBDBDBDB),
    .INIT_19(256'hE0E0E0E0E0E0E0E0E0DFDFDFDFDFDFDFDFDFDFDFDEDEDEDEDEDEDEDEDEDEDEDD),
    .INIT_1A(256'hE3E3E3E3E3E3E3E2E2E2E2E2E2E2E2E2E2E2E1E1E1E1E1E1E1E1E1E1E1E0E0E0),
    .INIT_1B(256'hE6E6E6E6E6E6E5E5E5E5E5E5E5E5E5E5E5E4E4E4E4E4E4E4E4E4E4E4E3E3E3E3),
    .INIT_1C(256'hE9E9E9E9E9E8E8E8E8E8E8E8E8E8E8E8E7E7E7E7E7E7E7E7E7E7E7E6E6E6E6E6),
    .INIT_1D(256'hECECECECEBEBEBEBEBEBEBEBEBEBEBEAEAEAEAEAEAEAEAEAEAEAE9E9E9E9E9E9),
    .INIT_1E(256'hEFEFEFEEEEEEEEEEEEEEEEEEEEEEEDEDEDEDEDEDEDEDEDEDEDECECECECECECEC),
    .INIT_1F(256'hF2F2F1F1F1F1F1F1F1F1F1F1F1F0F0F0F0F0F0F0F0F0F0F0EFEFEFEFEFEFEFEF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_036864_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_Naddra_o_al_n68 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i36_008,inst_doa_i36_007,inst_doa_i36_006,inst_doa_i36_005,inst_doa_i36_004,inst_doa_i36_003,inst_doa_i36_002,inst_doa_i36_001,inst_doa_i36_000}));
  // address_offset=37888;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'hF5F5F4F4F4F4F4F4F4F4F4F4F4F3F3F3F3F3F3F3F3F3F3F3F2F2F2F2F2F2F2F2),
    .INIT_01(256'hF8F8F7F7F7F7F7F7F7F7F7F7F7F6F6F6F6F6F6F6F6F6F6F5F5F5F5F5F5F5F5F5),
    .INIT_02(256'hFBFBFAFAFAFAFAFAFAFAFAFAFAF9F9F9F9F9F9F9F9F9F9F8F8F8F8F8F8F8F8F8),
    .INIT_03(256'hFEFEFDFDFDFDFDFDFDFDFDFDFDFCFCFCFCFCFCFCFCFCFCFBFBFBFBFBFBFBFBFB),
    .INIT_04(256'h01010000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFEFEFEFEFEFEFEFE),
    .INIT_05(256'h0404040303030303030303030302020202020202020202020101010101010101),
    .INIT_06(256'h0707070706060606060606060606050505050505050505050504040404040404),
    .INIT_07(256'h0A0A0A0A0A090909090909090909090808080808080808080807070707070707),
    .INIT_08(256'h0D0D0D0D0D0D0C0C0C0C0C0C0C0C0C0C0B0B0B0B0B0B0B0B0B0B0A0A0A0A0A0A),
    .INIT_09(256'h101010101010100F0F0F0F0F0F0F0F0F0F0E0E0E0E0E0E0E0E0E0E0D0D0D0D0D),
    .INIT_0A(256'h1313131313131313121212121212121212121111111111111111111111101010),
    .INIT_0B(256'h1616161616161616161615151515151515151515141414141414141414141313),
    .INIT_0C(256'h1A19191919191919191919181818181818181818181817171717171717171717),
    .INIT_0D(256'h1D1D1D1C1C1C1C1C1C1C1C1C1C1B1B1B1B1B1B1B1B1B1B1A1A1A1A1A1A1A1A1A),
    .INIT_0E(256'h20202020201F1F1F1F1F1F1F1F1F1F1E1E1E1E1E1E1E1E1E1E1D1D1D1D1D1D1D),
    .INIT_0F(256'h2323232323232322222222222222222222212121212121212121212020202020),
    .INIT_10(256'h2626262626262626262625252525252525252525242424242424242424242323),
    .INIT_11(256'h2A2A292929292929292929292828282828282828282827272727272727272727),
    .INIT_12(256'h2D2D2D2D2D2C2C2C2C2C2C2C2C2C2C2B2B2B2B2B2B2B2B2B2B2A2A2A2A2A2A2A),
    .INIT_13(256'h30303030303030302F2F2F2F2F2F2F2F2F2E2E2E2E2E2E2E2E2E2E2D2D2D2D2D),
    .INIT_14(256'h3433333333333333333333323232323232323232313131313131313131313030),
    .INIT_15(256'h3737373736363636363636363636353535353535353535343434343434343434),
    .INIT_16(256'h3A3A3A3A3A3A3A39393939393939393939383838383838383838373737373737),
    .INIT_17(256'h3E3D3D3D3D3D3D3D3D3D3D3C3C3C3C3C3C3C3C3C3B3B3B3B3B3B3B3B3B3B3A3A),
    .INIT_18(256'h41414141414040404040404040403F3F3F3F3F3F3F3F3F3F3E3E3E3E3E3E3E3E),
    .INIT_19(256'h4444444444444444434343434343434343434242424242424242424141414141),
    .INIT_1A(256'h4848474747474747474747474646464646464646464545454545454545454544),
    .INIT_1B(256'h4B4B4B4B4B4B4A4A4A4A4A4A4A4A4A4A49494949494949494948484848484848),
    .INIT_1C(256'h4F4E4E4E4E4E4E4E4E4E4D4D4D4D4D4D4D4D4D4D4C4C4C4C4C4C4C4C4C4B4B4B),
    .INIT_1D(256'h5252525252515151515151515151505050505050505050504F4F4F4F4F4F4F4F),
    .INIT_1E(256'h5555555555555555555454545454545454545453535353535353535352525252),
    .INIT_1F(256'h5959595959585858585858585858575757575757575757565656565656565656),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_037888_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_Naddra_o_al_n68 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i37_008,inst_doa_i37_007,inst_doa_i37_006,inst_doa_i37_005,inst_doa_i37_004,inst_doa_i37_003,inst_doa_i37_002,inst_doa_i37_001,inst_doa_i37_000}));
  // address_offset=38912;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'h5C5C5C5C5C5C5C5C5C5B5B5B5B5B5B5B5B5B5A5A5A5A5A5A5A5A5A5A59595959),
    .INIT_01(256'h60606060605F5F5F5F5F5F5F5F5F5E5E5E5E5E5E5E5E5E5D5D5D5D5D5D5D5D5D),
    .INIT_02(256'h6363636363636363636362626262626262626261616161616161616160606060),
    .INIT_03(256'h6767676767666666666666666666656565656565656565646464646464646464),
    .INIT_04(256'h6B6A6A6A6A6A6A6A6A6A69696969696969696968686868686868686867676767),
    .INIT_05(256'h6E6E6E6E6E6E6E6D6D6D6D6D6D6D6D6D6C6C6C6C6C6C6C6C6B6B6B6B6B6B6B6B),
    .INIT_06(256'h7272727171717171717171717070707070707070706F6F6F6F6F6F6F6F6F6E6E),
    .INIT_07(256'h7575757575757575747474747474747474737373737373737373727272727272),
    .INIT_08(256'h7979797979787878787878787878777777777777777777767676767676767675),
    .INIT_09(256'h7D7D7C7C7C7C7C7C7C7C7C7B7B7B7B7B7B7B7B7A7A7A7A7A7A7A7A7A79797979),
    .INIT_0A(256'h80808080808080807F7F7F7F7F7F7F7F7E7E7E7E7E7E7E7E7E7D7D7D7D7D7D7D),
    .INIT_0B(256'h8484848484838383838383838382828282828282828281818181818181818180),
    .INIT_0C(256'h8888878787878787878787868686868686868685858585858585858584848484),
    .INIT_0D(256'h8B8B8B8B8B8B8B8B8A8A8A8A8A8A8A8A8A898989898989898988888888888888),
    .INIT_0E(256'h8F8F8F8F8F8F8E8E8E8E8E8E8E8E8D8D8D8D8D8D8D8D8D8C8C8C8C8C8C8C8C8B),
    .INIT_0F(256'h93939392929292929292929291919191919191919090909090909090908F8F8F),
    .INIT_10(256'h9796969696969696969695959595959595959494949494949494949393939393),
    .INIT_11(256'h9A9A9A9A9A9A9A9A999999999999999998989898989898989897979797979797),
    .INIT_12(256'h9E9E9E9E9E9E9D9D9D9D9D9D9D9D9C9C9C9C9C9C9C9C9C9B9B9B9B9B9B9B9B9A),
    .INIT_13(256'hA2A2A2A2A1A1A1A1A1A1A1A1A0A0A0A0A0A0A0A0A09F9F9F9F9F9F9F9F9E9E9E),
    .INIT_14(256'hA6A6A5A5A5A5A5A5A5A5A5A4A4A4A4A4A4A4A4A3A3A3A3A3A3A3A3A2A2A2A2A2),
    .INIT_15(256'hAAA9A9A9A9A9A9A9A9A8A8A8A8A8A8A8A8A8A7A7A7A7A7A7A7A7A6A6A6A6A6A6),
    .INIT_16(256'hADADADADADADADADACACACACACACACACABABABABABABABABABAAAAAAAAAAAAAA),
    .INIT_17(256'hB1B1B1B1B1B1B1B0B0B0B0B0B0B0B0AFAFAFAFAFAFAFAFAEAEAEAEAEAEAEAEAE),
    .INIT_18(256'hB5B5B5B5B5B5B4B4B4B4B4B4B4B4B3B3B3B3B3B3B3B3B2B2B2B2B2B2B2B2B1B1),
    .INIT_19(256'hB9B9B9B9B9B8B8B8B8B8B8B8B8B7B7B7B7B7B7B7B7B6B6B6B6B6B6B6B6B5B5B5),
    .INIT_1A(256'hBDBDBDBDBCBCBCBCBCBCBCBCBBBBBBBBBBBBBBBBBABABABABABABABAB9B9B9B9),
    .INIT_1B(256'hC1C1C1C0C0C0C0C0C0C0C0BFBFBFBFBFBFBFBFBEBEBEBEBEBEBEBEBEBDBDBDBD),
    .INIT_1C(256'hC5C5C5C4C4C4C4C4C4C4C4C3C3C3C3C3C3C3C3C2C2C2C2C2C2C2C2C1C1C1C1C1),
    .INIT_1D(256'hC9C9C8C8C8C8C8C8C8C8C7C7C7C7C7C7C7C7C6C6C6C6C6C6C6C6C5C5C5C5C5C5),
    .INIT_1E(256'hCDCDCCCCCCCCCCCCCCCCCBCBCBCBCBCBCBCBCACACACACACACACAC9C9C9C9C9C9),
    .INIT_1F(256'hD1D1D0D0D0D0D0D0D0D0CFCFCFCFCFCFCFCFCECECECECECECECECDCDCDCDCDCD),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_038912_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_Naddra_o_al_n68 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i38_008,inst_doa_i38_007,inst_doa_i38_006,inst_doa_i38_005,inst_doa_i38_004,inst_doa_i38_003,inst_doa_i38_002,inst_doa_i38_001,inst_doa_i38_000}));
  // address_offset=39936;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'h000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hD5D5D4D4D4D4D4D4D4D4D3D3D3D3D3D3D3D3D2D2D2D2D2D2D2D2D1D1D1D1D1D1),
    .INIT_01(256'hD9D9D8D8D8D8D8D8D8D8D7D7D7D7D7D7D7D7D6D6D6D6D6D6D6D6D5D5D5D5D5D5),
    .INIT_02(256'hDDDDDCDCDCDCDCDCDCDCDBDBDBDBDBDBDBDBDADADADADADADADAD9D9D9D9D9D9),
    .INIT_03(256'hE1E1E0E0E0E0E0E0E0E0DFDFDFDFDFDFDFDFDEDEDEDEDEDEDEDEDDDDDDDDDDDD),
    .INIT_04(256'hE5E5E4E4E4E4E4E4E4E4E3E3E3E3E3E3E3E3E2E2E2E2E2E2E2E2E1E1E1E1E1E1),
    .INIT_05(256'hE9E9E9E8E8E8E8E8E8E8E8E7E7E7E7E7E7E7E7E6E6E6E6E6E6E6E6E5E5E5E5E5),
    .INIT_06(256'hEDEDEDEDECECECECECECECEBEBEBEBEBEBEBEBEAEAEAEAEAEAEAEAE9E9E9E9E9),
    .INIT_07(256'hF1F1F1F1F0F0F0F0F0F0F0F0EFEFEFEFEFEFEFEFEEEEEEEEEEEEEEEEEDEDEDED),
    .INIT_08(256'hF5F5F5F5F5F4F4F4F4F4F4F4F4F3F3F3F3F3F3F3F3F2F2F2F2F2F2F2F1F1F1F1),
    .INIT_09(256'hF9F9F9F9F9F9F8F8F8F8F8F8F8F8F7F7F7F7F7F7F7F7F6F6F6F6F6F6F6F5F5F5),
    .INIT_0A(256'hFDFDFDFDFDFDFDFCFCFCFCFCFCFCFCFBFBFBFBFBFBFBFBFAFAFAFAFAFAFAF9F9),
    .INIT_0B(256'h02010101010101010000000000000000FFFFFFFFFFFFFFFFFEFEFEFEFEFEFEFD),
    .INIT_0C(256'h0606050505050505050504040404040404030303030303030302020202020202),
    .INIT_0D(256'h0A0A0A0909090909090909080808080808080807070707070707060606060606),
    .INIT_0E(256'h0E0E0E0E0E0D0D0D0D0D0D0D0C0C0C0C0C0C0C0C0B0B0B0B0B0B0B0B0A0A0A0A),
    .INIT_0F(256'h121212121212111111111111111110101010101010100F0F0F0F0F0F0F0E0E0E),
    .INIT_10(256'h1616161616161616151515151515151514141414141414131313131313131312),
    .INIT_11(256'h1B1B1A1A1A1A1A1A1A1A19191919191919181818181818181817171717171717),
    .INIT_12(256'h1F1F1F1F1E1E1E1E1E1E1E1E1D1D1D1D1D1D1D1C1C1C1C1C1C1C1C1B1B1B1B1B),
    .INIT_13(256'h23232323232322222222222222222121212121212120202020202020201F1F1F),
    .INIT_14(256'h2827272727272727262626262626262625252525252525242424242424242423),
    .INIT_15(256'h2C2C2C2B2B2B2B2B2B2B2A2A2A2A2A2A2A2A2929292929292928282828282828),
    .INIT_16(256'h30303030302F2F2F2F2F2F2F2F2E2E2E2E2E2E2E2D2D2D2D2D2D2D2D2C2C2C2C),
    .INIT_17(256'h3434343434343434333333333333333232323232323231313131313131313030),
    .INIT_18(256'h3939393838383838383837373737373737373636363636363635353535353535),
    .INIT_19(256'h3D3D3D3D3D3C3C3C3C3C3C3C3C3B3B3B3B3B3B3B3A3A3A3A3A3A3A3939393939),
    .INIT_1A(256'h4241414141414141404040404040403F3F3F3F3F3F3F3F3E3E3E3E3E3E3E3D3D),
    .INIT_1B(256'h4646464545454545454545444444444444444343434343434342424242424242),
    .INIT_1C(256'h4A4A4A4A4A4A4949494949494949484848484848484747474747474746464646),
    .INIT_1D(256'h4F4F4E4E4E4E4E4E4E4D4D4D4D4D4D4D4C4C4C4C4C4C4C4C4B4B4B4B4B4B4B4A),
    .INIT_1E(256'h5353535353525252525252525151515151515150505050505050504F4F4F4F4F),
    .INIT_1F(256'h5857575757575757565656565656565555555555555555545454545454545353),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_039936_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_Naddra_o_al_n68 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i39_008,inst_doa_i39_007,inst_doa_i39_006,inst_doa_i39_005,inst_doa_i39_004,inst_doa_i39_003,inst_doa_i39_002,inst_doa_i39_001,inst_doa_i39_000}));
  // address_offset=40960;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h5C5C5C5C5B5B5B5B5B5B5B5A5A5A5A5A5A5A5A59595959595959585858585858),
    .INIT_01(256'h606060606060605F5F5F5F5F5F5F5F5E5E5E5E5E5E5E5D5D5D5D5D5D5D5C5C5C),
    .INIT_02(256'h6565656564646464646464636363636363636262626262626261616161616161),
    .INIT_03(256'h6969696969696968686868686868676767676767676666666666666666656565),
    .INIT_04(256'h6E6E6E6E6D6D6D6D6D6D6D6C6C6C6C6C6C6C6B6B6B6B6B6B6B6A6A6A6A6A6A6A),
    .INIT_05(256'h7272727272727271717171717171707070707070706F6F6F6F6F6F6F6F6E6E6E),
    .INIT_06(256'h7777777776767676767676757575757575757474747474747473737373737373),
    .INIT_07(256'h7C7B7B7B7B7B7B7B7A7A7A7A7A7A7A7979797979797978787878787878777777),
    .INIT_08(256'h80808080807F7F7F7F7F7F7F7E7E7E7E7E7E7E7D7D7D7D7D7D7D7C7C7C7C7C7C),
    .INIT_09(256'h8585848484848484848383838383838382828282828282818181818181818080),
    .INIT_0A(256'h8989898989898888888888888887878787878787868686868686868585858585),
    .INIT_0B(256'h8E8E8E8D8D8D8D8D8D8D8C8C8C8C8C8C8C8B8B8B8B8B8B8B8A8A8A8A8A8A8A89),
    .INIT_0C(256'h9292929292929291919191919191909090909090908F8F8F8F8F8F8F8E8E8E8E),
    .INIT_0D(256'h9797979796969696969696959595959595959494949494949493939393939393),
    .INIT_0E(256'h9C9C9B9B9B9B9B9B9B9A9A9A9A9A9A9A99999999999999989898989898979797),
    .INIT_0F(256'hA0A0A0A0A0A09F9F9F9F9F9F9F9E9E9E9E9E9E9E9D9D9D9D9D9D9D9C9C9C9C9C),
    .INIT_10(256'hA5A5A5A5A4A4A4A4A4A4A4A3A3A3A3A3A3A3A2A2A2A2A2A2A2A1A1A1A1A1A1A0),
    .INIT_11(256'hAAAAA9A9A9A9A9A9A9A8A8A8A8A8A8A7A7A7A7A7A7A7A6A6A6A6A6A6A6A5A5A5),
    .INIT_12(256'hAEAEAEAEAEAEADADADADADADADACACACACACACACABABABABABABABAAAAAAAAAA),
    .INIT_13(256'hB3B3B3B3B2B2B2B2B2B2B2B1B1B1B1B1B1B1B0B0B0B0B0B0B0AFAFAFAFAFAFAF),
    .INIT_14(256'hB8B8B7B7B7B7B7B7B7B6B6B6B6B6B6B6B5B5B5B5B5B5B5B4B4B4B4B4B4B3B3B3),
    .INIT_15(256'hBCBCBCBCBCBCBCBBBBBBBBBBBBBBBABABABABABABAB9B9B9B9B9B9B9B8B8B8B8),
    .INIT_16(256'hC1C1C1C1C1C0C0C0C0C0C0C0BFBFBFBFBFBFBFBEBEBEBEBEBEBEBDBDBDBDBDBD),
    .INIT_17(256'hC6C6C6C6C5C5C5C5C5C5C4C4C4C4C4C4C4C3C3C3C3C3C3C3C2C2C2C2C2C2C2C1),
    .INIT_18(256'hCBCBCACACACACACACAC9C9C9C9C9C9C9C8C8C8C8C8C8C7C7C7C7C7C7C7C6C6C6),
    .INIT_19(256'hD0CFCFCFCFCFCFCECECECECECECECDCDCDCDCDCDCDCCCCCCCCCCCCCBCBCBCBCB),
    .INIT_1A(256'hD4D4D4D4D4D4D3D3D3D3D3D3D3D2D2D2D2D2D2D1D1D1D1D1D1D1D0D0D0D0D0D0),
    .INIT_1B(256'hD9D9D9D9D9D8D8D8D8D8D8D7D7D7D7D7D7D7D6D6D6D6D6D6D6D5D5D5D5D5D5D4),
    .INIT_1C(256'hDEDEDEDDDDDDDDDDDDDDDCDCDCDCDCDCDCDBDBDBDBDBDBDADADADADADADAD9D9),
    .INIT_1D(256'hE3E3E2E2E2E2E2E2E2E1E1E1E1E1E1E0E0E0E0E0E0E0DFDFDFDFDFDFDFDEDEDE),
    .INIT_1E(256'hE8E7E7E7E7E7E7E7E6E6E6E6E6E6E5E5E5E5E5E5E5E4E4E4E4E4E4E3E3E3E3E3),
    .INIT_1F(256'hECECECECECECECEBEBEBEBEBEBEAEAEAEAEAEAEAE9E9E9E9E9E9E8E8E8E8E8E8),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_040960_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_addra_o_al_n76 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i40_008,inst_doa_i40_007,inst_doa_i40_006,inst_doa_i40_005,inst_doa_i40_004,inst_doa_i40_003,inst_doa_i40_002,inst_doa_i40_001,inst_doa_i40_000}));
  // address_offset=40960;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'h0000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_040960_009 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n2484,open_n2485,open_n2486,open_n2487,open_n2488,open_n2489,open_n2490,1'b0,open_n2491}),
    .rsta(rsta),
    .doa({open_n2506,open_n2507,open_n2508,open_n2509,open_n2510,open_n2511,open_n2512,open_n2513,inst_doa_i40_009}));
  // address_offset=40960;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000000000000000000),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_040960_010 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n2542,open_n2543,open_n2544,open_n2545,open_n2546,open_n2547,open_n2548,1'b0,open_n2549}),
    .rsta(rsta),
    .doa({open_n2564,open_n2565,open_n2566,open_n2567,open_n2568,open_n2569,open_n2570,open_n2571,inst_doa_i40_010}));
  // address_offset=40960;data_offset=11;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_040960_011 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n2600,open_n2601,open_n2602,open_n2603,open_n2604,open_n2605,open_n2606,1'b0,open_n2607}),
    .rsta(rsta),
    .doa({open_n2622,open_n2623,open_n2624,open_n2625,open_n2626,open_n2627,open_n2628,open_n2629,inst_doa_i40_011}));
  // address_offset=41984;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000000000000000),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'hF1F1F1F1F1F1F0F0F0F0F0F0EFEFEFEFEFEFEFEEEEEEEEEEEEEDEDEDEDEDEDED),
    .INIT_01(256'hF6F6F6F6F6F5F5F5F5F5F5F4F4F4F4F4F4F4F3F3F3F3F3F3F3F2F2F2F2F2F2F1),
    .INIT_02(256'hFBFBFBFBFAFAFAFAFAFAFAF9F9F9F9F9F9F8F8F8F8F8F8F8F7F7F7F7F7F7F6F6),
    .INIT_03(256'h000000FFFFFFFFFFFFFFFEFEFEFEFEFEFDFDFDFDFDFDFDFCFCFCFCFCFCFCFBFB),
    .INIT_04(256'h0505050404040404040303030303030302020202020201010101010101000000),
    .INIT_05(256'h0A0A090909090909090808080808080707070707070706060606060605050505),
    .INIT_06(256'h0F0F0E0E0E0E0E0E0D0D0D0D0D0D0D0C0C0C0C0C0C0B0B0B0B0B0B0B0A0A0A0A),
    .INIT_07(256'h1414131313131313121212121212111111111111111010101010100F0F0F0F0F),
    .INIT_08(256'h1918181818181818171717171717161616161616161515151515151414141414),
    .INIT_09(256'h1E1D1D1D1D1D1D1C1C1C1C1C1C1C1B1B1B1B1B1B1A1A1A1A1A1A1A1919191919),
    .INIT_0A(256'h23222222222222212121212121212020202020201F1F1F1F1F1F1F1E1E1E1E1E),
    .INIT_0B(256'h2827272727272726262626262626252525252525242424242424242323232323),
    .INIT_0C(256'h2D2C2C2C2C2C2C2B2B2B2B2B2B2B2A2A2A2A2A2A292929292929282828282828),
    .INIT_0D(256'h32313131313131303030303030302F2F2F2F2F2F2E2E2E2E2E2E2E2D2D2D2D2D),
    .INIT_0E(256'h3736363636363636353535353535343434343434333333333333333232323232),
    .INIT_0F(256'h3C3B3B3B3B3B3B3B3A3A3A3A3A3A393939393939383838383838383737373737),
    .INIT_10(256'h41414040404040403F3F3F3F3F3F3E3E3E3E3E3E3E3D3D3D3D3D3D3C3C3C3C3C),
    .INIT_11(256'h4646454545454545444444444444444343434343434242424242424141414141),
    .INIT_12(256'h4B4B4B4A4A4A4A4A4A4949494949494848484848484847474747474746464646),
    .INIT_13(256'h5050504F4F4F4F4F4F4E4E4E4E4E4E4E4D4D4D4D4D4D4C4C4C4C4C4C4B4B4B4B),
    .INIT_14(256'h5555555554545454545453535353535352525252525252515151515151505050),
    .INIT_15(256'h5A5A5A5A59595959595959585858585858575757575757565656565656555555),
    .INIT_16(256'h5F5F5F5F5F5E5E5E5E5E5E5D5D5D5D5D5D5D5C5C5C5C5C5C5B5B5B5B5B5B5A5A),
    .INIT_17(256'h646464646464636363636363626262626262616161616161616060606060605F),
    .INIT_18(256'h6A69696969696968686868686867676767676766666666666665656565656565),
    .INIT_19(256'h6F6F6E6E6E6E6E6E6D6D6D6D6D6D6C6C6C6C6C6C6B6B6B6B6B6B6A6A6A6A6A6A),
    .INIT_1A(256'h7474747373737373737272727272727171717171717070707070706F6F6F6F6F),
    .INIT_1B(256'h7979797978787878787877777777777776767676767675757575757574747474),
    .INIT_1C(256'h7E7E7E7E7E7D7D7D7D7D7D7C7C7C7C7C7C7B7B7B7B7B7B7A7A7A7A7A7A797979),
    .INIT_1D(256'h8383838383838282828282828181818181818080808080807F7F7F7F7F7F7F7E),
    .INIT_1E(256'h8988888888888887878787878786868686868685858585858585848484848484),
    .INIT_1F(256'h8E8E8D8D8D8D8D8D8D8C8C8C8C8C8C8B8B8B8B8B8B8A8A8A8A8A8A8989898989),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_041984_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_addra_o_al_n76 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i41_008,inst_doa_i41_007,inst_doa_i41_006,inst_doa_i41_005,inst_doa_i41_004,inst_doa_i41_003,inst_doa_i41_002,inst_doa_i41_001,inst_doa_i41_000}));
  // address_offset=43008;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'h0000000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h939393939292929292929191919191919090909090908F8F8F8F8F8F8E8E8E8E),
    .INIT_01(256'h9898989898979797979797969696969696959595959595959494949494949393),
    .INIT_02(256'h9E9D9D9D9D9D9D9C9C9C9C9C9C9B9B9B9B9B9B9A9A9A9A9A9A99999999999998),
    .INIT_03(256'hA3A3A2A2A2A2A2A2A1A1A1A1A1A1A0A0A0A0A0A09F9F9F9F9F9F9F9E9E9E9E9E),
    .INIT_04(256'hA8A8A8A8A7A7A7A7A7A7A6A6A6A6A6A6A5A5A5A5A5A5A4A4A4A4A4A4A3A3A3A3),
    .INIT_05(256'hADADADADADADACACACACACACABABABABABABAAAAAAAAAAAAA9A9A9A9A9A9A8A8),
    .INIT_06(256'hB3B2B2B2B2B2B2B1B1B1B1B1B1B0B0B0B0B0B0AFAFAFAFAFAFAEAEAEAEAEAEAD),
    .INIT_07(256'hB8B8B8B7B7B7B7B7B7B6B6B6B6B6B6B5B5B5B5B5B5B4B4B4B4B4B4B3B3B3B3B3),
    .INIT_08(256'hBDBDBDBDBDBCBCBCBCBCBCBBBBBBBBBBBBBABABABABABAB9B9B9B9B9B9B8B8B8),
    .INIT_09(256'hC3C2C2C2C2C2C2C1C1C1C1C1C1C0C0C0C0C0C0BFBFBFBFBFBFBEBEBEBEBEBEBD),
    .INIT_0A(256'hC8C8C8C7C7C7C7C7C7C6C6C6C6C6C6C5C5C5C5C5C5C4C4C4C4C4C4C3C3C3C3C3),
    .INIT_0B(256'hCDCDCDCDCDCCCCCCCCCCCCCBCBCBCBCBCBCACACACACACAC9C9C9C9C9C9C8C8C8),
    .INIT_0C(256'hD3D2D2D2D2D2D2D1D1D1D1D1D1D0D0D0D0D0D0CFCFCFCFCFCFCECECECECECECD),
    .INIT_0D(256'hD8D8D8D7D7D7D7D7D7D6D6D6D6D6D6D5D5D5D5D5D5D4D4D4D4D4D4D3D3D3D3D3),
    .INIT_0E(256'hDDDDDDDDDDDCDCDCDCDCDCDBDBDBDBDBDBDADADADADADAD9D9D9D9D9D9D8D8D8),
    .INIT_0F(256'hE3E3E2E2E2E2E2E2E1E1E1E1E1E1E0E0E0E0E0E0DFDFDFDFDFDFDEDEDEDEDEDD),
    .INIT_10(256'hE8E8E8E8E7E7E7E7E7E7E6E6E6E6E6E6E5E5E5E5E5E5E4E4E4E4E4E4E3E3E3E3),
    .INIT_11(256'hEEEDEDEDEDEDECECECECECECEBEBEBEBEBEBEAEAEAEAEAEAE9E9E9E9E9E9E8E8),
    .INIT_12(256'hF3F3F3F2F2F2F2F2F2F1F1F1F1F1F1F0F0F0F0F0F0EFEFEFEFEFEFEEEEEEEEEE),
    .INIT_13(256'hF8F8F8F8F8F7F7F7F7F7F7F6F6F6F6F6F6F5F5F5F5F5F5F4F4F4F4F4F4F3F3F3),
    .INIT_14(256'hFEFEFDFDFDFDFDFDFCFCFCFCFCFCFBFBFBFBFBFBFAFAFAFAFAFAF9F9F9F9F9F9),
    .INIT_15(256'h03030303030202020202020101010101000000000000FFFFFFFFFFFFFEFEFEFE),
    .INIT_16(256'h0908080808080807070707070706060606060605050505050504040404040403),
    .INIT_17(256'h0E0E0E0E0D0D0D0D0D0D0C0C0C0C0C0C0B0B0B0B0B0B0A0A0A0A0A0A09090909),
    .INIT_18(256'h1413131313131312121212121211111111111110101010100F0F0F0F0F0F0E0E),
    .INIT_19(256'h1919191918181818181817171717171716161616161515151515151414141414),
    .INIT_1A(256'h1F1E1E1E1E1E1E1D1D1D1D1D1C1C1C1C1C1C1B1B1B1B1B1B1A1A1A1A1A1A1919),
    .INIT_1B(256'h2424242423232323232322222222222121212121212020202020201F1F1F1F1F),
    .INIT_1C(256'h2A29292929292928282828282727272727272626262626262525252525252424),
    .INIT_1D(256'h2F2F2F2F2E2E2E2E2E2E2D2D2D2D2D2C2C2C2C2C2C2B2B2B2B2B2B2A2A2A2A2A),
    .INIT_1E(256'h3534343434343433333333333332323232323131313131313030303030302F2F),
    .INIT_1F(256'h3A3A3A3A39393939393938383838383837373737373736363636363535353535),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_043008_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_addra_o_al_n76 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i42_008,inst_doa_i42_007,inst_doa_i42_006,inst_doa_i42_005,inst_doa_i42_004,inst_doa_i42_003,inst_doa_i42_002,inst_doa_i42_001,inst_doa_i42_000}));
  // address_offset=44032;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h40403F3F3F3F3F3E3E3E3E3E3E3D3D3D3D3D3D3C3C3C3C3C3C3B3B3B3B3B3A3A),
    .INIT_01(256'h4545454545444444444444434343434342424242424241414141414140404040),
    .INIT_02(256'h4B4B4A4A4A4A4A4A494949494949484848484847474747474746464646464645),
    .INIT_03(256'h5050505050504F4F4F4F4F4E4E4E4E4E4E4D4D4D4D4D4D4C4C4C4C4C4B4B4B4B),
    .INIT_04(256'h5656565555555555555454545454545353535353525252525252515151515151),
    .INIT_05(256'h5C5B5B5B5B5B5A5A5A5A5A5A5959595959595858585858585757575757565656),
    .INIT_06(256'h616161616060606060605F5F5F5F5F5F5E5E5E5E5E5D5D5D5D5D5D5C5C5C5C5C),
    .INIT_07(256'h6767666666666666656565656564646464646463636363636362626262626161),
    .INIT_08(256'h6C6C6C6C6C6B6B6B6B6B6B6A6A6A6A6A6A696969696968686868686867676767),
    .INIT_09(256'h7272727171717171717070707070706F6F6F6F6F6E6E6E6E6E6E6D6D6D6D6D6D),
    .INIT_0A(256'h7877777777777776767676767675757575757474747474747373737373737272),
    .INIT_0B(256'h7D7D7D7D7D7C7C7C7C7C7B7B7B7B7B7B7A7A7A7A7A7A79797979797878787878),
    .INIT_0C(256'h83838382828282828181818181818080808080807F7F7F7F7F7E7E7E7E7E7E7D),
    .INIT_0D(256'h8988888888888887878787878686868686868585858585848484848484838383),
    .INIT_0E(256'h8E8E8E8E8E8D8D8D8D8D8C8C8C8C8C8C8B8B8B8B8B8B8A8A8A8A8A8989898989),
    .INIT_0F(256'h949494939393939392929292929291919191919190909090908F8F8F8F8F8F8E),
    .INIT_10(256'h9A99999999999998989898989797979797979696969696969595959595949494),
    .INIT_11(256'h9F9F9F9F9F9E9E9E9E9E9D9D9D9D9D9D9C9C9C9C9C9C9B9B9B9B9B9A9A9A9A9A),
    .INIT_12(256'hA5A5A5A4A4A4A4A4A4A3A3A3A3A3A2A2A2A2A2A2A1A1A1A1A1A1A0A0A0A0A09F),
    .INIT_13(256'hABABAAAAAAAAAAA9A9A9A9A9A9A8A8A8A8A8A7A7A7A7A7A7A6A6A6A6A6A6A5A5),
    .INIT_14(256'hB0B0B0B0B0B0AFAFAFAFAFAEAEAEAEAEAEADADADADADACACACACACACABABABAB),
    .INIT_15(256'hB6B6B6B6B5B5B5B5B5B5B4B4B4B4B4B3B3B3B3B3B3B2B2B2B2B2B1B1B1B1B1B1),
    .INIT_16(256'hBCBCBBBBBBBBBBBBBABABABABABAB9B9B9B9B9B8B8B8B8B8B8B7B7B7B7B7B6B6),
    .INIT_17(256'hC2C1C1C1C1C1C1C0C0C0C0C0BFBFBFBFBFBFBEBEBEBEBEBDBDBDBDBDBDBCBCBC),
    .INIT_18(256'hC7C7C7C7C7C6C6C6C6C6C6C5C5C5C5C5C4C4C4C4C4C4C3C3C3C3C3C2C2C2C2C2),
    .INIT_19(256'hCDCDCDCDCCCCCCCCCCCBCBCBCBCBCBCACACACACAC9C9C9C9C9C9C8C8C8C8C8C8),
    .INIT_1A(256'hD3D3D2D2D2D2D2D2D1D1D1D1D1D1D0D0D0D0D0CFCFCFCFCFCFCECECECECECDCD),
    .INIT_1B(256'hD9D8D8D8D8D8D8D7D7D7D7D7D6D6D6D6D6D6D5D5D5D5D5D4D4D4D4D4D4D3D3D3),
    .INIT_1C(256'hDEDEDEDEDEDDDDDDDDDDDDDCDCDCDCDCDCDBDBDBDBDBDADADADADADAD9D9D9D9),
    .INIT_1D(256'hE4E4E4E4E3E3E3E3E3E3E2E2E2E2E2E1E1E1E1E1E1E0E0E0E0E0DFDFDFDFDFDF),
    .INIT_1E(256'hEAEAEAE9E9E9E9E9E9E8E8E8E8E8E7E7E7E7E7E7E6E6E6E6E6E5E5E5E5E5E5E4),
    .INIT_1F(256'hF0F0EFEFEFEFEFEFEEEEEEEEEEEDEDEDEDEDEDECECECECECEBEBEBEBEBEBEAEA),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_044032_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_addra_o_al_n76 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i43_008,inst_doa_i43_007,inst_doa_i43_006,inst_doa_i43_005,inst_doa_i43_004,inst_doa_i43_003,inst_doa_i43_002,inst_doa_i43_001,inst_doa_i43_000}));
  // address_offset=45056;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'hF6F5F5F5F5F5F4F4F4F4F4F4F3F3F3F3F3F2F2F2F2F2F2F1F1F1F1F1F0F0F0F0),
    .INIT_01(256'hFBFBFBFBFBFAFAFAFAFAFAF9F9F9F9F9F8F8F8F8F8F8F7F7F7F7F7F6F6F6F6F6),
    .INIT_02(256'h01010101000000000000FFFFFFFFFFFEFEFEFEFEFEFDFDFDFDFDFCFCFCFCFCFC),
    .INIT_03(256'h0707070606060606060505050505040404040404030303030302020202020201),
    .INIT_04(256'h0D0D0D0C0C0C0C0C0B0B0B0B0B0B0A0A0A0A0A09090909090908080808080707),
    .INIT_05(256'h1313121212121211111111111110101010100F0F0F0F0F0F0E0E0E0E0E0D0D0D),
    .INIT_06(256'h1918181818181717171717171616161616151515151515141414141413131313),
    .INIT_07(256'h1E1E1E1E1E1E1D1D1D1D1D1C1C1C1C1C1C1B1B1B1B1B1A1A1A1A1A1919191919),
    .INIT_08(256'h2424242424232323232322222222222221212121212020202020201F1F1F1F1F),
    .INIT_09(256'h2A2A2A2A29292929292928282828282727272727262626262626252525252524),
    .INIT_0A(256'h3030302F2F2F2F2F2F2E2E2E2E2E2D2D2D2D2D2D2C2C2C2C2C2B2B2B2B2B2B2A),
    .INIT_0B(256'h3636363535353535343434343434333333333332323232323231313131313030),
    .INIT_0C(256'h3C3C3B3B3B3B3B3B3A3A3A3A3A39393939393938383838383737373737363636),
    .INIT_0D(256'h424241414141414040404040403F3F3F3F3F3E3E3E3E3E3D3D3D3D3D3D3C3C3C),
    .INIT_0E(256'h4847474747474746464646464545454545444444444444434343434342424242),
    .INIT_0F(256'h4E4D4D4D4D4D4C4C4C4C4C4C4B4B4B4B4B4A4A4A4A4A49494949494948484848),
    .INIT_10(256'h535353535353525252525251515151515050505050504F4F4F4F4F4E4E4E4E4E),
    .INIT_11(256'h5959595959585858585858575757575756565656565555555555555454545454),
    .INIT_12(256'h5F5F5F5F5F5E5E5E5E5E5D5D5D5D5D5D5C5C5C5C5C5B5B5B5B5B5A5A5A5A5A5A),
    .INIT_13(256'h656565656464646464646363636363626262626262616161616160606060605F),
    .INIT_14(256'h6B6B6B6B6A6A6A6A6A6A69696969696868686868676767676767666666666665),
    .INIT_15(256'h7171717170707070706F6F6F6F6F6F6E6E6E6E6E6D6D6D6D6D6C6C6C6C6C6C6B),
    .INIT_16(256'h7777777776767676767575757575747474747474737373737372727272727271),
    .INIT_17(256'h7D7D7D7C7C7C7C7C7C7B7B7B7B7B7A7A7A7A7A7A797979797978787878787777),
    .INIT_18(256'h838383828282828282818181818180808080807F7F7F7F7F7F7E7E7E7E7E7D7D),
    .INIT_19(256'h8989898888888888878787878787868686868685858585858584848484848383),
    .INIT_1A(256'h8F8F8F8E8E8E8E8E8D8D8D8D8D8D8C8C8C8C8C8B8B8B8B8B8A8A8A8A8A8A8989),
    .INIT_1B(256'h9595959494949494939393939393929292929291919191919090909090908F8F),
    .INIT_1C(256'h9B9B9B9A9A9A9A9A999999999999989898989897979797979696969696969595),
    .INIT_1D(256'hA1A1A1A0A0A0A0A09F9F9F9F9F9F9E9E9E9E9E9D9D9D9D9D9C9C9C9C9C9C9B9B),
    .INIT_1E(256'hA7A7A7A6A6A6A6A6A5A5A5A5A5A5A4A4A4A4A4A3A3A3A3A3A2A2A2A2A2A2A1A1),
    .INIT_1F(256'hADADADACACACACACABABABABABABAAAAAAAAAAA9A9A9A9A9A8A8A8A8A8A8A7A7),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_045056_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_addra[_o_al_n84 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i44_008,inst_doa_i44_007,inst_doa_i44_006,inst_doa_i44_005,inst_doa_i44_004,inst_doa_i44_003,inst_doa_i44_002,inst_doa_i44_001,inst_doa_i44_000}));
  // address_offset=46080;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'h0000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hB3B3B3B2B2B2B2B2B1B1B1B1B1B1B0B0B0B0B0AFAFAFAFAFAEAEAEAEAEAEADAD),
    .INIT_01(256'hB9B9B9B8B8B8B8B8B7B7B7B7B7B7B6B6B6B6B6B5B5B5B5B5B4B4B4B4B4B4B3B3),
    .INIT_02(256'hBFBFBFBEBEBEBEBEBEBDBDBDBDBDBCBCBCBCBCBBBBBBBBBBBABABABABABAB9B9),
    .INIT_03(256'hC5C5C5C4C4C4C4C4C4C3C3C3C3C3C2C2C2C2C2C1C1C1C1C1C1C0C0C0C0C0BFBF),
    .INIT_04(256'hCBCBCBCBCACACACACAC9C9C9C9C9C8C8C8C8C8C7C7C7C7C7C7C6C6C6C6C6C5C5),
    .INIT_05(256'hD1D1D1D1D0D0D0D0D0CFCFCFCFCFCECECECECECECDCDCDCDCDCCCCCCCCCCCBCB),
    .INIT_06(256'hD7D7D7D7D6D6D6D6D6D5D5D5D5D5D5D4D4D4D4D4D3D3D3D3D3D2D2D2D2D2D1D1),
    .INIT_07(256'hDDDDDDDDDCDCDCDCDCDCDBDBDBDBDBDADADADADAD9D9D9D9D9D8D8D8D8D8D8D7),
    .INIT_08(256'hE3E3E3E3E3E2E2E2E2E2E1E1E1E1E1E0E0E0E0E0DFDFDFDFDFDFDEDEDEDEDEDD),
    .INIT_09(256'hE9E9E9E9E9E8E8E8E8E8E7E7E7E7E7E6E6E6E6E6E6E5E5E5E5E5E4E4E4E4E4E3),
    .INIT_0A(256'hEFEFEFEFEFEEEEEEEEEEEEEDEDEDEDEDECECECECECEBEBEBEBEBEAEAEAEAEAEA),
    .INIT_0B(256'hF5F5F5F5F5F5F4F4F4F4F4F3F3F3F3F3F2F2F2F2F2F1F1F1F1F1F1F0F0F0F0F0),
    .INIT_0C(256'hFCFBFBFBFBFBFAFAFAFAFAF9F9F9F9F9F9F8F8F8F8F8F7F7F7F7F7F6F6F6F6F6),
    .INIT_0D(256'h020101010101000000000000FFFFFFFFFFFEFEFEFEFEFDFDFDFDFDFCFCFCFCFC),
    .INIT_0E(256'h0808070707070706060606060505050505040404040404030303030302020202),
    .INIT_0F(256'h0E0E0D0D0D0D0D0C0C0C0C0C0C0B0B0B0B0B0A0A0A0A0A090909090908080808),
    .INIT_10(256'h1414141313131313121212121211111111111010101010100F0F0F0F0F0E0E0E),
    .INIT_11(256'h1A1A1A1919191919181818181818171717171716161616161515151515141414),
    .INIT_12(256'h202020201F1F1F1F1F1E1E1E1E1E1D1D1D1D1D1C1C1C1C1C1C1B1B1B1B1B1A1A),
    .INIT_13(256'h2626262625252525252424242424242323232323222222222221212121212020),
    .INIT_14(256'h2C2C2C2C2C2B2B2B2B2B2A2A2A2A2A2929292929292828282828272727272726),
    .INIT_15(256'h323232323231313131313130303030302F2F2F2F2F2E2E2E2E2E2D2D2D2D2D2D),
    .INIT_16(256'h3938383838383737373737363636363636353535353534343434343333333333),
    .INIT_17(256'h3F3F3E3E3E3E3E3D3D3D3D3D3C3C3C3C3C3B3B3B3B3B3A3A3A3A3A3A39393939),
    .INIT_18(256'h454544444444444343434343434242424242414141414140404040403F3F3F3F),
    .INIT_19(256'h4B4B4B4A4A4A4A4A494949494948484848484847474747474646464646454545),
    .INIT_1A(256'h5151515150505050504F4F4F4F4F4E4E4E4E4E4D4D4D4D4D4C4C4C4C4C4C4B4B),
    .INIT_1B(256'h5757575756565656565655555555555454545454535353535352525252525151),
    .INIT_1C(256'h5D5D5D5D5D5C5C5C5C5C5B5B5B5B5B5B5A5A5A5A5A5959595959585858585857),
    .INIT_1D(256'h646363636363626262626261616161616060606060605F5F5F5F5F5E5E5E5E5E),
    .INIT_1E(256'h6A6A696969696968686868686767676767666666666665656565656564646464),
    .INIT_1F(256'h70706F6F6F6F6F6F6E6E6E6E6E6D6D6D6D6D6C6C6C6C6C6B6B6B6B6B6A6A6A6A),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_046080_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_addra[_o_al_n84 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i45_008,inst_doa_i45_007,inst_doa_i45_006,inst_doa_i45_005,inst_doa_i45_004,inst_doa_i45_003,inst_doa_i45_002,inst_doa_i45_001,inst_doa_i45_000}));
  // address_offset=47104;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'hFFFFFFE000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'h7676767575757575747474747474737373737372727272727171717171707070),
    .INIT_01(256'h7C7C7C7C7B7B7B7B7B7A7A7A7A7A797979797979787878787877777777777676),
    .INIT_02(256'h8282828282818181818180808080807F7F7F7F7F7F7E7E7E7E7E7D7D7D7D7D7C),
    .INIT_03(256'h8988888888888787878787868686868685858585858484848484848383838383),
    .INIT_04(256'h8F8F8E8E8E8E8E8D8D8D8D8D8C8C8C8C8C8B8B8B8B8B8A8A8A8A8A8989898989),
    .INIT_05(256'h959595949494949493939393939292929292919191919190909090908F8F8F8F),
    .INIT_06(256'h9B9B9B9A9A9A9A9A9A9999999999989898989897979797979696969696959595),
    .INIT_07(256'hA1A1A1A1A0A0A0A0A0A09F9F9F9F9F9E9E9E9E9E9D9D9D9D9D9C9C9C9C9C9B9B),
    .INIT_08(256'hA7A7A7A7A7A6A6A6A6A6A6A5A5A5A5A5A4A4A4A4A4A3A3A3A3A3A2A2A2A2A2A1),
    .INIT_09(256'hAEADADADADADACACACACACACABABABABABAAAAAAAAAAA9A9A9A9A9A8A8A8A8A8),
    .INIT_0A(256'hB4B4B3B3B3B3B3B2B2B2B2B2B2B1B1B1B1B1B0B0B0B0B0AFAFAFAFAFAEAEAEAE),
    .INIT_0B(256'hBABABAB9B9B9B9B9B8B8B8B8B8B8B7B7B7B7B7B6B6B6B6B6B5B5B5B5B5B4B4B4),
    .INIT_0C(256'hC0C0C0C0BFBFBFBFBFBFBEBEBEBEBEBDBDBDBDBDBCBCBCBCBCBBBBBBBBBBBABA),
    .INIT_0D(256'hC6C6C6C6C6C5C5C5C5C5C5C4C4C4C4C4C3C3C3C3C3C2C2C2C2C2C1C1C1C1C1C0),
    .INIT_0E(256'hCDCCCCCCCCCCCBCBCBCBCBCBCACACACACAC9C9C9C9C9C8C8C8C8C8C7C7C7C7C7),
    .INIT_0F(256'hD3D3D2D2D2D2D2D2D1D1D1D1D1D0D0D0D0D0CFCFCFCFCFCECECECECECDCDCDCD),
    .INIT_10(256'hD9D9D9D9D8D8D8D8D8D7D7D7D7D7D6D6D6D6D6D5D5D5D5D5D4D4D4D4D4D3D3D3),
    .INIT_11(256'hDFDFDFDFDFDEDEDEDEDEDDDDDDDDDDDCDCDCDCDCDBDBDBDBDBDADADADADAD9D9),
    .INIT_12(256'hE6E5E5E5E5E5E4E4E4E4E4E3E3E3E3E3E2E2E2E2E2E1E1E1E1E1E0E0E0E0E0E0),
    .INIT_13(256'hECECEBEBEBEBEBEAEAEAEAEAE9E9E9E9E9E8E8E8E8E8E7E7E7E7E7E7E6E6E6E6),
    .INIT_14(256'hF2F2F2F1F1F1F1F1F0F0F0F0F0EFEFEFEFEFEEEEEEEEEEEEEDEDEDEDEDECECEC),
    .INIT_15(256'hF8F8F8F8F7F7F7F7F7F6F6F6F6F6F5F5F5F5F5F5F4F4F4F4F4F3F3F3F3F3F2F2),
    .INIT_16(256'hFEFEFEFEFEFDFDFDFDFDFCFCFCFCFCFCFBFBFBFBFBFAFAFAFAFAF9F9F9F9F9F8),
    .INIT_17(256'h050404040404040303030303020202020201010101010000000000FFFFFFFFFF),
    .INIT_18(256'h0B0B0B0A0A0A0A0A090909090908080808080707070707060606060605050505),
    .INIT_19(256'h1111111110101010100F0F0F0F0F0E0E0E0E0E0D0D0D0D0D0C0C0C0C0C0B0B0B),
    .INIT_1A(256'h1717171717161616161615151515151414141414131313131313121212121211),
    .INIT_1B(256'h1E1D1D1D1D1D1C1C1C1C1C1B1B1B1B1B1B1A1A1A1A1A19191919191818181818),
    .INIT_1C(256'h24242323232323232222222222212121212120202020201F1F1F1F1F1E1E1E1E),
    .INIT_1D(256'h2A2A2A2A29292929292828282828272727272726262626262525252525242424),
    .INIT_1E(256'h30303030302F2F2F2F2F2E2E2E2E2E2D2D2D2D2D2C2C2C2C2C2B2B2B2B2B2B2A),
    .INIT_1F(256'h3736363636363535353535343434343433333333333332323232323131313131),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_047104_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_addra[_o_al_n84 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i46_008,inst_doa_i46_007,inst_doa_i46_006,inst_doa_i46_005,inst_doa_i46_004,inst_doa_i46_003,inst_doa_i46_002,inst_doa_i46_001,inst_doa_i46_000}));
  // address_offset=48128;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'h3D3D3C3C3C3C3C3B3B3B3B3B3B3A3A3A3A3A3939393939383838383837373737),
    .INIT_01(256'h434343434242424242414141414140404040403F3F3F3F3F3E3E3E3E3E3D3D3D),
    .INIT_02(256'h4949494949484848484847474747474646464646454545454544444444444443),
    .INIT_03(256'h504F4F4F4F4F4E4E4E4E4E4D4D4D4D4D4D4C4C4C4C4C4B4B4B4B4B4A4A4A4A4A),
    .INIT_04(256'h5656565555555555545454545453535353535252525252515151515150505050),
    .INIT_05(256'h5C5C5C5C5B5B5B5B5B5A5A5A5A5A595959595958585858585757575757565656),
    .INIT_06(256'h6262626262616161616160606060605F5F5F5F5F5F5E5E5E5E5E5D5D5D5D5D5C),
    .INIT_07(256'h6968686868686867676767676666666666656565656564646464646363636363),
    .INIT_08(256'h6F6F6F6E6E6E6E6E6D6D6D6D6D6C6C6C6C6C6B6B6B6B6B6A6A6A6A6A69696969),
    .INIT_09(256'h7575757574747474747373737373727272727271717171717170707070706F6F),
    .INIT_0A(256'h7B7B7B7B7B7B7A7A7A7A7A797979797978787878787777777777767676767675),
    .INIT_0B(256'h8282818181818180808080807F7F7F7F7F7E7E7E7E7E7D7D7D7D7D7C7C7C7C7C),
    .INIT_0C(256'h8888888787878787868686868685858585858484848484848383838383828282),
    .INIT_0D(256'h8E8E8E8E8E8D8D8D8D8D8C8C8C8C8C8B8B8B8B8B8A8A8A8A8A89898989898888),
    .INIT_0E(256'h95949494949493939393939292929292919191919190909090908F8F8F8F8F8E),
    .INIT_0F(256'h9B9B9A9A9A9A9A99999999999898989898989797979797969696969695959595),
    .INIT_10(256'hA1A1A1A1A0A0A0A0A09F9F9F9F9F9E9E9E9E9E9D9D9D9D9D9C9C9C9C9C9B9B9B),
    .INIT_11(256'hA7A7A7A7A7A6A6A6A6A6A5A5A5A5A5A4A4A4A4A4A3A3A3A3A3A2A2A2A2A2A2A1),
    .INIT_12(256'hAEADADADADADACACACACACACABABABABABAAAAAAAAAAA9A9A9A9A9A8A8A8A8A8),
    .INIT_13(256'hB4B4B4B3B3B3B3B3B2B2B2B2B2B1B1B1B1B1B0B0B0B0B0AFAFAFAFAFAEAEAEAE),
    .INIT_14(256'hBABABABAB9B9B9B9B9B8B8B8B8B8B7B7B7B7B7B6B6B6B6B6B6B5B5B5B5B5B4B4),
    .INIT_15(256'hC0C0C0C0C0C0BFBFBFBFBFBEBEBEBEBEBDBDBDBDBDBCBCBCBCBCBBBBBBBBBBBA),
    .INIT_16(256'hC7C7C6C6C6C6C6C5C5C5C5C5C4C4C4C4C4C3C3C3C3C3C2C2C2C2C2C1C1C1C1C1),
    .INIT_17(256'hCDCDCDCCCCCCCCCCCBCBCBCBCBCBCACACACACAC9C9C9C9C9C8C8C8C8C8C7C7C7),
    .INIT_18(256'hD3D3D3D3D3D2D2D2D2D2D1D1D1D1D1D0D0D0D0D0CFCFCFCFCFCECECECECECDCD),
    .INIT_19(256'hDAD9D9D9D9D9D8D8D8D8D8D7D7D7D7D7D6D6D6D6D6D5D5D5D5D5D5D4D4D4D4D4),
    .INIT_1A(256'hE0E0E0DFDFDFDFDFDEDEDEDEDEDDDDDDDDDDDCDCDCDCDCDBDBDBDBDBDADADADA),
    .INIT_1B(256'hE6E6E6E6E5E5E5E5E5E4E4E4E4E4E3E3E3E3E3E2E2E2E2E2E1E1E1E1E1E0E0E0),
    .INIT_1C(256'hECECECECECEBEBEBEBEBEAEAEAEAEAEAE9E9E9E9E9E8E8E8E8E8E7E7E7E7E7E6),
    .INIT_1D(256'hF3F3F2F2F2F2F2F1F1F1F1F1F0F0F0F0F0EFEFEFEFEFEEEEEEEEEEEDEDEDEDED),
    .INIT_1E(256'hF9F9F9F8F8F8F8F8F7F7F7F7F7F6F6F6F6F6F5F5F5F5F5F5F4F4F4F4F4F3F3F3),
    .INIT_1F(256'hFFFFFFFFFFFEFEFEFEFEFDFDFDFDFDFCFCFCFCFCFBFBFBFBFBFAFAFAFAFAF9F9),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_048128_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_addra[_o_al_n84 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i47_008,inst_doa_i47_007,inst_doa_i47_006,inst_doa_i47_005,inst_doa_i47_004,inst_doa_i47_003,inst_doa_i47_002,inst_doa_i47_001,inst_doa_i47_000}));
  // address_offset=49152;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0605050505050404040404030303030302020202020101010101000000000000),
    .INIT_01(256'h0C0C0B0B0B0B0B0A0A0A0A0A0A09090909090808080808070707070706060606),
    .INIT_02(256'h12121212111111111110101010100F0F0F0F0F0E0E0E0E0E0D0D0D0D0D0C0C0C),
    .INIT_03(256'h1818181818171717171716161616161515151515151414141414131313131312),
    .INIT_04(256'h1F1F1E1E1E1E1E1D1D1D1D1D1C1C1C1C1C1B1B1B1B1B1A1A1A1A1A1919191919),
    .INIT_05(256'h252525242424242423232323232222222222212121212120202020201F1F1F1F),
    .INIT_06(256'h2B2B2B2B2A2A2A2A2A2A29292929292828282828272727272726262626262525),
    .INIT_07(256'h32313131313130303030302F2F2F2F2F2E2E2E2E2E2D2D2D2D2D2C2C2C2C2C2B),
    .INIT_08(256'h3838373737373736363636363535353535343434343434333333333332323232),
    .INIT_09(256'h3E3E3E3E3D3D3D3D3D3C3C3C3C3C3B3B3B3B3B3A3A3A3A3A3939393939383838),
    .INIT_0A(256'h444444444443434343434242424242414141414140404040403F3F3F3F3F3F3E),
    .INIT_0B(256'h4B4A4A4A4A4A4949494949494848484848474747474746464646464545454545),
    .INIT_0C(256'h51515150505050504F4F4F4F4F4E4E4E4E4E4D4D4D4D4D4C4C4C4C4C4B4B4B4B),
    .INIT_0D(256'h5757575756565656565555555555545454545453535353535352525252525151),
    .INIT_0E(256'h5D5D5D5D5D5D5C5C5C5C5C5B5B5B5B5B5A5A5A5A5A5959595959585858585857),
    .INIT_0F(256'h646463636363636262626262616161616160606060605F5F5F5F5F5E5E5E5E5E),
    .INIT_10(256'h6A6A6A6969696969686868686867676767676766666666666565656565646464),
    .INIT_11(256'h70707070706F6F6F6F6F6E6E6E6E6E6D6D6D6D6D6C6C6C6C6C6B6B6B6B6B6A6A),
    .INIT_12(256'h7776767676767575757575747474747473737373737272727272717171717171),
    .INIT_13(256'h7D7D7C7C7C7C7C7B7B7B7B7B7B7A7A7A7A7A7979797979787878787877777777),
    .INIT_14(256'h838383838282828282818181818180808080807F7F7F7F7F7E7E7E7E7E7D7D7D),
    .INIT_15(256'h8989898989888888888887878787878686868686858585858584848484848483),
    .INIT_16(256'h908F8F8F8F8F8E8E8E8E8E8E8D8D8D8D8D8C8C8C8C8C8B8B8B8B8B8A8A8A8A8A),
    .INIT_17(256'h9696969595959595949494949493939393939292929292919191919190909090),
    .INIT_18(256'h9C9C9C9C9B9B9B9B9B9A9A9A9A9A999999999998989898989797979797979696),
    .INIT_19(256'hA2A2A2A2A2A1A1A1A1A1A0A0A0A0A0A09F9F9F9F9F9E9E9E9E9E9D9D9D9D9D9C),
    .INIT_1A(256'hA9A9A8A8A8A8A8A7A7A7A7A7A6A6A6A6A6A5A5A5A5A5A4A4A4A4A4A3A3A3A3A3),
    .INIT_1B(256'hAFAFAFAEAEAEAEAEADADADADADACACACACACABABABABABAAAAAAAAAAA9A9A9A9),
    .INIT_1C(256'hB5B5B5B5B4B4B4B4B4B3B3B3B3B3B2B2B2B2B2B2B1B1B1B1B1B0B0B0B0B0AFAF),
    .INIT_1D(256'hBBBBBBBBBBBBBABABABABAB9B9B9B9B9B8B8B8B8B8B7B7B7B7B7B6B6B6B6B6B5),
    .INIT_1E(256'hC2C2C1C1C1C1C1C0C0C0C0C0BFBFBFBFBFBEBEBEBEBEBDBDBDBDBDBCBCBCBCBC),
    .INIT_1F(256'hC8C8C8C7C7C7C7C7C6C6C6C6C6C5C5C5C5C5C4C4C4C4C4C4C3C3C3C3C3C2C2C2),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_049152_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_Naddr_o_al_n92 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i48_008,inst_doa_i48_007,inst_doa_i48_006,inst_doa_i48_005,inst_doa_i48_004,inst_doa_i48_003,inst_doa_i48_002,inst_doa_i48_001,inst_doa_i48_000}));
  // address_offset=49152;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000000000000),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'h0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_049152_009 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n2994,open_n2995,open_n2996,open_n2997,open_n2998,open_n2999,open_n3000,1'b0,open_n3001}),
    .rsta(rsta),
    .doa({open_n3016,open_n3017,open_n3018,open_n3019,open_n3020,open_n3021,open_n3022,open_n3023,inst_doa_i48_009}));
  // address_offset=49152;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000000000000000000000),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_049152_010 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n3052,open_n3053,open_n3054,open_n3055,open_n3056,open_n3057,open_n3058,1'b0,open_n3059}),
    .rsta(rsta),
    .doa({open_n3074,open_n3075,open_n3076,open_n3077,open_n3078,open_n3079,open_n3080,open_n3081,inst_doa_i48_010}));
  // address_offset=49152;data_offset=11;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_049152_011 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n3110,open_n3111,open_n3112,open_n3113,open_n3114,open_n3115,open_n3116,1'b0,open_n3117}),
    .rsta(rsta),
    .doa({open_n3132,open_n3133,open_n3134,open_n3135,open_n3136,open_n3137,open_n3138,open_n3139,inst_doa_i48_011}));
  // address_offset=50176;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'hCECECECECDCDCDCDCDCCCCCCCCCCCCCBCBCBCBCBCACACACACAC9C9C9C9C9C8C8),
    .INIT_01(256'hD4D4D4D4D4D4D3D3D3D3D3D2D2D2D2D2D1D1D1D1D1D0D0D0D0D0CFCFCFCFCFCE),
    .INIT_02(256'hDBDBDADADADADAD9D9D9D9D9D8D8D8D8D8D7D7D7D7D7D6D6D6D6D6D5D5D5D5D5),
    .INIT_03(256'hE1E1E1E0E0E0E0E0DFDFDFDFDFDEDEDEDEDEDDDDDDDDDDDCDCDCDCDCDCDBDBDB),
    .INIT_04(256'hE7E7E7E7E6E6E6E6E6E5E5E5E5E5E4E4E4E4E4E4E3E3E3E3E3E2E2E2E2E2E1E1),
    .INIT_05(256'hEDEDEDEDEDECECECECECECEBEBEBEBEBEAEAEAEAEAE9E9E9E9E9E8E8E8E8E8E7),
    .INIT_06(256'hF4F4F3F3F3F3F3F2F2F2F2F2F1F1F1F1F1F0F0F0F0F0EFEFEFEFEFEEEEEEEEEE),
    .INIT_07(256'hFAFAFAF9F9F9F9F9F8F8F8F8F8F7F7F7F7F7F6F6F6F6F6F5F5F5F5F5F4F4F4F4),
    .INIT_08(256'h00000000FFFFFFFFFFFEFEFEFEFEFDFDFDFDFDFCFCFCFCFCFBFBFBFBFBFBFAFA),
    .INIT_09(256'h0606060606050505050504040404040303030303030202020202010101010100),
    .INIT_0A(256'h0D0C0C0C0C0C0B0B0B0B0B0A0A0A0A0A0A090909090908080808080707070707),
    .INIT_0B(256'h1313121212121211111111111110101010100F0F0F0F0F0E0E0E0E0E0D0D0D0D),
    .INIT_0C(256'h1919191818181818181717171717161616161615151515151414141414131313),
    .INIT_0D(256'h1F1F1F1F1F1E1E1E1E1E1D1D1D1D1D1C1C1C1C1C1B1B1B1B1B1A1A1A1A1A1919),
    .INIT_0E(256'h262525252525242424242423232323232222222222212121212120202020201F),
    .INIT_0F(256'h2C2C2B2B2B2B2B2A2A2A2A2A2929292929282828282827272727272626262626),
    .INIT_10(256'h323232313131313130303030302F2F2F2F2F2E2E2E2E2E2D2D2D2D2D2D2C2C2C),
    .INIT_11(256'h3838383837373737373636363636353535353534343434343433333333333232),
    .INIT_12(256'h3E3E3E3E3E3D3D3D3D3D3C3C3C3C3C3B3B3B3B3B3A3A3A3A3A3A393939393938),
    .INIT_13(256'h4544444444444343434343424242424241414141414040404040403F3F3F3F3F),
    .INIT_14(256'h4B4B4A4A4A4A4A49494949494848484848474747474747464646464645454545),
    .INIT_15(256'h51515150505050504F4F4F4F4F4E4E4E4E4E4D4D4D4D4D4D4C4C4C4C4C4B4B4B),
    .INIT_16(256'h5757575756565656565555555555545454545453535353535352525252525151),
    .INIT_17(256'h5D5D5D5D5D5C5C5C5C5C5B5B5B5B5B5A5A5A5A5A595959595959585858585857),
    .INIT_18(256'h6463636363636262626262616161616160606060605F5F5F5F5F5F5E5E5E5E5E),
    .INIT_19(256'h6A6A696969696968686868686767676767666666666665656565656564646464),
    .INIT_1A(256'h7070706F6F6F6F6F6E6E6E6E6E6D6D6D6D6D6C6C6C6C6C6B6B6B6B6B6A6A6A6A),
    .INIT_1B(256'h7676767675757575757474747474737373737372727272727171717171707070),
    .INIT_1C(256'h7C7C7C7C7B7B7B7B7B7B7A7A7A7A7A7979797979787878787877777777777676),
    .INIT_1D(256'h828282828281818181818080808080807F7F7F7F7F7E7E7E7E7E7D7D7D7D7D7C),
    .INIT_1E(256'h8988888888888787878787868686868686858585858584848484848383838383),
    .INIT_1F(256'h8F8F8E8E8E8E8E8D8D8D8D8D8C8C8C8C8C8B8B8B8B8B8B8A8A8A8A8A89898989),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_050176_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_Naddr_o_al_n92 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i49_008,inst_doa_i49_007,inst_doa_i49_006,inst_doa_i49_005,inst_doa_i49_004,inst_doa_i49_003,inst_doa_i49_002,inst_doa_i49_001,inst_doa_i49_000}));
  // address_offset=51200;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'h000000000000000000000000000000000000000000001FFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h95959594949494949393939393929292929291919191919090909090908F8F8F),
    .INIT_01(256'h9B9B9B9A9A9A9A9A9A9999999999989898989897979797979696969696959595),
    .INIT_02(256'hA1A1A1A1A0A0A0A0A09F9F9F9F9F9F9E9E9E9E9E9D9D9D9D9D9C9C9C9C9C9B9B),
    .INIT_03(256'hA7A7A7A7A7A6A6A6A6A6A5A5A5A5A5A4A4A4A4A4A4A3A3A3A3A3A2A2A2A2A2A1),
    .INIT_04(256'hAEADADADADADACACACACACABABABABABAAAAAAAAAAA9A9A9A9A9A9A8A8A8A8A8),
    .INIT_05(256'hB4B3B3B3B3B3B3B2B2B2B2B2B1B1B1B1B1B0B0B0B0B0AFAFAFAFAFAEAEAEAEAE),
    .INIT_06(256'hBABAB9B9B9B9B9B8B8B8B8B8B7B7B7B7B7B7B6B6B6B6B6B5B5B5B5B5B4B4B4B4),
    .INIT_07(256'hC0C0C0BFBFBFBFBFBEBEBEBEBEBDBDBDBDBDBCBCBCBCBCBCBBBBBBBBBBBABABA),
    .INIT_08(256'hC6C6C6C5C5C5C5C5C5C4C4C4C4C4C3C3C3C3C3C2C2C2C2C2C1C1C1C1C1C0C0C0),
    .INIT_09(256'hCCCCCCCCCBCBCBCBCBCACACACACAC9C9C9C9C9C9C8C8C8C8C8C7C7C7C7C7C6C6),
    .INIT_0A(256'hD2D2D2D2D2D1D1D1D1D1D0D0D0D0D0CFCFCFCFCFCECECECECECECDCDCDCDCDCC),
    .INIT_0B(256'hD8D8D8D8D8D7D7D7D7D7D6D6D6D6D6D6D5D5D5D5D5D4D4D4D4D4D3D3D3D3D3D2),
    .INIT_0C(256'hDFDEDEDEDEDEDDDDDDDDDDDCDCDCDCDCDBDBDBDBDBDBDADADADADAD9D9D9D9D9),
    .INIT_0D(256'hE5E4E4E4E4E4E3E3E3E3E3E3E2E2E2E2E2E1E1E1E1E1E0E0E0E0E0DFDFDFDFDF),
    .INIT_0E(256'hEBEBEAEAEAEAEAE9E9E9E9E9E8E8E8E8E8E7E7E7E7E7E7E6E6E6E6E6E5E5E5E5),
    .INIT_0F(256'hF1F1F0F0F0F0F0EFEFEFEFEFEFEEEEEEEEEEEDEDEDEDEDECECECECECEBEBEBEB),
    .INIT_10(256'hF7F7F7F6F6F6F6F6F5F5F5F5F5F4F4F4F4F4F3F3F3F3F3F3F2F2F2F2F2F1F1F1),
    .INIT_11(256'hFDFDFDFCFCFCFCFCFBFBFBFBFBFBFAFAFAFAFAF9F9F9F9F9F8F8F8F8F8F7F7F7),
    .INIT_12(256'h03030303020202020201010101010000000000FFFFFFFFFFFFFEFEFEFEFEFDFD),
    .INIT_13(256'h0909090908080808080707070707060606060606050505050504040404040303),
    .INIT_14(256'h0F0F0F0F0E0E0E0E0E0E0D0D0D0D0D0C0C0C0C0C0B0B0B0B0B0A0A0A0A0A0A09),
    .INIT_15(256'h151515151514141414141313131313121212121211111111111110101010100F),
    .INIT_16(256'h1B1B1B1B1B1A1A1A1A1A19191919191918181818181717171717161616161615),
    .INIT_17(256'h21212121212020202020201F1F1F1F1F1E1E1E1E1E1D1D1D1D1D1C1C1C1C1C1C),
    .INIT_18(256'h2727272727272626262626252525252524242424242323232323232222222222),
    .INIT_19(256'h2E2D2D2D2D2D2C2C2C2C2C2B2B2B2B2B2A2A2A2A2A2A29292929292828282828),
    .INIT_1A(256'h343333333333323232323231313131313130303030302F2F2F2F2F2E2E2E2E2E),
    .INIT_1B(256'h3A39393939393838383838383737373737363636363635353535353434343434),
    .INIT_1C(256'h403F3F3F3F3F3E3E3E3E3E3E3D3D3D3D3D3C3C3C3C3C3B3B3B3B3B3B3A3A3A3A),
    .INIT_1D(256'h4645454545454544444444444343434343424242424241414141414140404040),
    .INIT_1E(256'h4C4B4B4B4B4B4B4A4A4A4A4A4949494949484848484848474747474746464646),
    .INIT_1F(256'h5251515151515150505050504F4F4F4F4F4E4E4E4E4E4E4D4D4D4D4D4C4C4C4C),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_051200_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_Naddr_o_al_n92 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i50_008,inst_doa_i50_007,inst_doa_i50_006,inst_doa_i50_005,inst_doa_i50_004,inst_doa_i50_003,inst_doa_i50_002,inst_doa_i50_001,inst_doa_i50_000}));
  // address_offset=52224;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFF8000000000000000000000000000000000000000000),
    .INIT_00(256'h5857575757575756565656565555555555545454545454535353535352525252),
    .INIT_01(256'h5E5D5D5D5D5D5D5C5C5C5C5C5B5B5B5B5B5A5A5A5A5A5A595959595958585858),
    .INIT_02(256'h64636363636363626262626261616161616060606060605F5F5F5F5F5E5E5E5E),
    .INIT_03(256'h6A69696969696968686868686767676767666666666666656565656564646464),
    .INIT_04(256'h706F6F6F6F6F6F6E6E6E6E6E6D6D6D6D6D6C6C6C6C6C6C6B6B6B6B6B6A6A6A6A),
    .INIT_05(256'h7675757575757574747474747373737373727272727272717171717170707070),
    .INIT_06(256'h7C7B7B7B7B7B7A7A7A7A7A7A7979797979787878787878777777777776767676),
    .INIT_07(256'h8281818181818080808080807F7F7F7F7F7E7E7E7E7E7D7D7D7D7D7D7C7C7C7C),
    .INIT_08(256'h8887878787878686868686858585858585848484848483838383838382828282),
    .INIT_09(256'h8D8D8D8D8D8D8C8C8C8C8C8B8B8B8B8B8B8A8A8A8A8A89898989898888888888),
    .INIT_0A(256'h939393939393929292929291919191919090909090908F8F8F8F8F8E8E8E8E8E),
    .INIT_0B(256'h9999999999989898989898979797979796969696969595959595959494949494),
    .INIT_0C(256'h9F9F9F9F9F9E9E9E9E9E9D9D9D9D9D9D9C9C9C9C9C9B9B9B9B9B9B9A9A9A9A9A),
    .INIT_0D(256'hA5A5A5A5A5A4A4A4A4A4A3A3A3A3A3A2A2A2A2A2A2A1A1A1A1A1A0A0A0A0A0A0),
    .INIT_0E(256'hABABABABAAAAAAAAAAAAA9A9A9A9A9A8A8A8A8A8A7A7A7A7A7A7A6A6A6A6A6A5),
    .INIT_0F(256'hB1B1B1B1B0B0B0B0B0AFAFAFAFAFAFAEAEAEAEAEADADADADADACACACACACACAB),
    .INIT_10(256'hB7B7B7B6B6B6B6B6B6B5B5B5B5B5B4B4B4B4B4B3B3B3B3B3B3B2B2B2B2B2B1B1),
    .INIT_11(256'hBDBDBDBCBCBCBCBCBBBBBBBBBBBBBABABABABAB9B9B9B9B9B8B8B8B8B8B8B7B7),
    .INIT_12(256'hC3C3C2C2C2C2C2C2C1C1C1C1C1C0C0C0C0C0BFBFBFBFBFBFBEBEBEBEBEBDBDBD),
    .INIT_13(256'hC9C9C8C8C8C8C8C7C7C7C7C7C6C6C6C6C6C6C5C5C5C5C5C4C4C4C4C4C4C3C3C3),
    .INIT_14(256'hCFCECECECECECDCDCDCDCDCDCCCCCCCCCCCBCBCBCBCBCBCACACACACAC9C9C9C9),
    .INIT_15(256'hD4D4D4D4D4D4D3D3D3D3D3D2D2D2D2D2D2D1D1D1D1D1D0D0D0D0D0D0CFCFCFCF),
    .INIT_16(256'hDADADADADAD9D9D9D9D9D9D8D8D8D8D8D7D7D7D7D7D6D6D6D6D6D6D5D5D5D5D5),
    .INIT_17(256'hE0E0E0E0DFDFDFDFDFDFDEDEDEDEDEDDDDDDDDDDDDDCDCDCDCDCDBDBDBDBDBDB),
    .INIT_18(256'hE6E6E6E6E5E5E5E5E5E4E4E4E4E4E3E3E3E3E3E3E2E2E2E2E2E1E1E1E1E1E1E0),
    .INIT_19(256'hECECECEBEBEBEBEBEAEAEAEAEAEAE9E9E9E9E9E8E8E8E8E8E8E7E7E7E7E7E6E6),
    .INIT_1A(256'hF2F2F1F1F1F1F1F0F0F0F0F0F0EFEFEFEFEFEEEEEEEEEEEEEDEDEDEDEDECECEC),
    .INIT_1B(256'hF8F7F7F7F7F7F6F6F6F6F6F6F5F5F5F5F5F4F4F4F4F4F4F3F3F3F3F3F2F2F2F2),
    .INIT_1C(256'hFDFDFDFDFDFDFCFCFCFCFCFBFBFBFBFBFBFAFAFAFAFAF9F9F9F9F9F9F8F8F8F8),
    .INIT_1D(256'h030303030302020202020101010101010000000000FFFFFFFFFFFFFEFEFEFEFE),
    .INIT_1E(256'h0909090908080808080707070707070606060606050505050505040404040403),
    .INIT_1F(256'h0F0F0F0E0E0E0E0E0D0D0D0D0D0D0C0C0C0C0C0B0B0B0B0B0B0A0A0A0A0A0909),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_052224_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_Naddr_o_al_n92 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i51_008,inst_doa_i51_007,inst_doa_i51_006,inst_doa_i51_005,inst_doa_i51_004,inst_doa_i51_003,inst_doa_i51_002,inst_doa_i51_001,inst_doa_i51_000}));
  // address_offset=53248;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'h15141414141414131313131312121212121211111111111010101010100F0F0F),
    .INIT_01(256'h1A1A1A1A1A1A1919191919181818181818171717171716161616161615151515),
    .INIT_02(256'h20202020201F1F1F1F1F1E1E1E1E1E1E1D1D1D1D1D1C1C1C1C1C1C1B1B1B1B1B),
    .INIT_03(256'h2626262525252525252424242424232323232323222222222222212121212120),
    .INIT_04(256'h2C2C2B2B2B2B2B2B2A2A2A2A2A29292929292928282828282727272727272626),
    .INIT_05(256'h3231313131313030303030302F2F2F2F2F2E2E2E2E2E2E2D2D2D2D2D2D2C2C2C),
    .INIT_06(256'h3737373737363636363636353535353534343434343433333333333232323232),
    .INIT_07(256'h3D3D3D3D3C3C3C3C3C3B3B3B3B3B3B3A3A3A3A3A393939393939383838383837),
    .INIT_08(256'h434342424242424241414141414040404040403F3F3F3F3F3E3E3E3E3E3E3D3D),
    .INIT_09(256'h4948484848484747474747474646464646454545454545444444444444434343),
    .INIT_0A(256'h4E4E4E4E4E4D4D4D4D4D4C4C4C4C4C4C4B4B4B4B4B4A4A4A4A4A4A4949494949),
    .INIT_0B(256'h545454535353535353525252525251515151515150505050504F4F4F4F4F4F4E),
    .INIT_0C(256'h5A59595959595958585858585857575757575656565656565555555555545454),
    .INIT_0D(256'h5F5F5F5F5F5E5E5E5E5E5E5D5D5D5D5D5D5C5C5C5C5C5B5B5B5B5B5B5A5A5A5A),
    .INIT_0E(256'h6565656564646464646363636363636262626262626161616161606060606060),
    .INIT_0F(256'h6B6B6A6A6A6A6A69696969696968686868686867676767676666666666666565),
    .INIT_10(256'h7070707070706F6F6F6F6F6E6E6E6E6E6E6D6D6D6D6D6D6C6C6C6C6C6B6B6B6B),
    .INIT_11(256'h7676767675757575757474747474747373737373737272727272717171717171),
    .INIT_12(256'h7C7C7B7B7B7B7B7B7A7A7A7A7A79797979797978787878787777777777777676),
    .INIT_13(256'h81818181818180808080807F7F7F7F7F7F7E7E7E7E7E7E7D7D7D7D7D7C7C7C7C),
    .INIT_14(256'h8787878786868686868585858585858484848484848383838383828282828282),
    .INIT_15(256'h8D8C8C8C8C8C8C8B8B8B8B8B8B8A8A8A8A8A8989898989898888888888888787),
    .INIT_16(256'h929292929291919191919190909090908F8F8F8F8F8F8E8E8E8E8E8E8D8D8D8D),
    .INIT_17(256'h9898989797979797979696969696959595959595949494949494939393939392),
    .INIT_18(256'h9E9D9D9D9D9D9C9C9C9C9C9C9B9B9B9B9B9B9A9A9A9A9A999999999999989898),
    .INIT_19(256'hA3A3A3A3A2A2A2A2A2A2A1A1A1A1A1A0A0A0A0A0A09F9F9F9F9F9F9E9E9E9E9E),
    .INIT_1A(256'hA9A9A8A8A8A8A8A7A7A7A7A7A7A6A6A6A6A6A6A5A5A5A5A5A5A4A4A4A4A4A3A3),
    .INIT_1B(256'hAEAEAEAEAEADADADADADADACACACACACABABABABABABAAAAAAAAAAAAA9A9A9A9),
    .INIT_1C(256'hB4B4B4B3B3B3B3B3B2B2B2B2B2B2B1B1B1B1B1B1B0B0B0B0B0AFAFAFAFAFAFAE),
    .INIT_1D(256'hB9B9B9B9B9B9B8B8B8B8B8B8B7B7B7B7B7B6B6B6B6B6B6B5B5B5B5B5B5B4B4B4),
    .INIT_1E(256'hBFBFBFBEBEBEBEBEBEBDBDBDBDBDBDBCBCBCBCBCBBBBBBBBBBBBBABABABABABA),
    .INIT_1F(256'hC5C4C4C4C4C4C3C3C3C3C3C3C2C2C2C2C2C2C1C1C1C1C1C1C0C0C0C0C0BFBFBF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_053248_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_Naddra_o_al_n100 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i52_008,inst_doa_i52_007,inst_doa_i52_006,inst_doa_i52_005,inst_doa_i52_004,inst_doa_i52_003,inst_doa_i52_002,inst_doa_i52_001,inst_doa_i52_000}));
  // address_offset=54272;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'h0000000000000000000000000000000000000000007FFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hCACACACAC9C9C9C9C9C8C8C8C8C8C8C7C7C7C7C7C7C6C6C6C6C6C6C5C5C5C5C5),
    .INIT_01(256'hD0CFCFCFCFCFCFCECECECECECECDCDCDCDCDCCCCCCCCCCCCCBCBCBCBCBCBCACA),
    .INIT_02(256'hD5D5D5D5D4D4D4D4D4D4D3D3D3D3D3D3D2D2D2D2D2D1D1D1D1D1D1D0D0D0D0D0),
    .INIT_03(256'hDBDADADADADADAD9D9D9D9D9D9D8D8D8D8D8D8D7D7D7D7D7D6D6D6D6D6D6D5D5),
    .INIT_04(256'hE0E0E0E0DFDFDFDFDFDFDEDEDEDEDEDEDDDDDDDDDDDCDCDCDCDCDCDBDBDBDBDB),
    .INIT_05(256'hE6E5E5E5E5E5E5E4E4E4E4E4E4E3E3E3E3E3E3E2E2E2E2E2E1E1E1E1E1E1E0E0),
    .INIT_06(256'hEBEBEBEBEAEAEAEAEAEAE9E9E9E9E9E9E8E8E8E8E8E7E7E7E7E7E7E6E6E6E6E6),
    .INIT_07(256'hF1F0F0F0F0F0F0EFEFEFEFEFEEEEEEEEEEEEEDEDEDEDEDEDECECECECECECEBEB),
    .INIT_08(256'hF6F6F6F5F5F5F5F5F5F4F4F4F4F4F4F3F3F3F3F3F3F2F2F2F2F2F2F1F1F1F1F1),
    .INIT_09(256'hFBFBFBFBFBFBFAFAFAFAFAFAF9F9F9F9F9F9F8F8F8F8F8F8F7F7F7F7F7F7F6F6),
    .INIT_0A(256'h010101000000000000FFFFFFFFFFFFFEFEFEFEFEFDFDFDFDFDFDFCFCFCFCFCFC),
    .INIT_0B(256'h0606060606050505050505040404040404030303030303020202020202010101),
    .INIT_0C(256'h0C0C0B0B0B0B0B0B0A0A0A0A0A0A090909090909080808080808070707070706),
    .INIT_0D(256'h111111111010101010100F0F0F0F0F0F0E0E0E0E0E0E0D0D0D0D0D0D0C0C0C0C),
    .INIT_0E(256'h1716161616161615151515151514141414141413131313131312121212121111),
    .INIT_0F(256'h1C1C1C1B1B1B1B1B1B1A1A1A1A1A1A1919191919191818181818181717171717),
    .INIT_10(256'h21212121212020202020201F1F1F1F1F1F1E1E1E1E1E1E1D1D1D1D1D1D1C1C1C),
    .INIT_11(256'h2727262626262626252525252525242424242424232323232323222222222222),
    .INIT_12(256'h2C2C2C2C2B2B2B2B2B2B2A2A2A2A2A2A29292929292928282828282827272727),
    .INIT_13(256'h3131313131313030303030302F2F2F2F2F2F2E2E2E2E2E2E2D2D2D2D2D2D2C2C),
    .INIT_14(256'h3737363636363636353535353535343434343434333333333333323232323232),
    .INIT_15(256'h3C3C3C3C3B3B3B3B3B3B3A3A3A3A3A3A39393939393938383838383837373737),
    .INIT_16(256'h4141414141414040404040403F3F3F3F3F3F3E3E3E3E3E3E3D3D3D3D3D3D3C3C),
    .INIT_17(256'h4747464646464646454545454545444444444444434343434343424242424242),
    .INIT_18(256'h4C4C4C4C4B4B4B4B4B4B4A4A4A4A4A4A49494949494948484848484847474747),
    .INIT_19(256'h5151515151515050505050504F4F4F4F4F4F4E4E4E4E4E4E4D4D4D4D4D4D4C4C),
    .INIT_1A(256'h5756565656565655555555555554545454545453535353535352525252525252),
    .INIT_1B(256'h5C5C5C5B5B5B5B5B5B5A5A5A5A5A5A5959595959595858585858585757575757),
    .INIT_1C(256'h61616161606060606060605F5F5F5F5F5F5E5E5E5E5E5E5D5D5D5D5D5D5C5C5C),
    .INIT_1D(256'h6666666666666565656565656464646464646363636363636262626262626161),
    .INIT_1E(256'h6C6B6B6B6B6B6B6A6A6A6A6A6A6A696969696969686868686868676767676767),
    .INIT_1F(256'h7171717070707070706F6F6F6F6F6F6E6E6E6E6E6E6D6D6D6D6D6D6C6C6C6C6C),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_054272_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_Naddra_o_al_n100 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i53_008,inst_doa_i53_007,inst_doa_i53_006,inst_doa_i53_005,inst_doa_i53_004,inst_doa_i53_003,inst_doa_i53_002,inst_doa_i53_001,inst_doa_i53_000}));
  // address_offset=55296;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000000000000),
    .INIT_00(256'h7676767675757575757574747474747473737373737372727272727272717171),
    .INIT_01(256'h7B7B7B7B7B7A7A7A7A7A7A7A7979797979797878787878787777777777777676),
    .INIT_02(256'h808080808080807F7F7F7F7F7F7E7E7E7E7E7E7D7D7D7D7D7D7C7C7C7C7C7C7B),
    .INIT_03(256'h8686858585858585848484848484838383838383828282828282818181818181),
    .INIT_04(256'h8B8B8B8A8A8A8A8A8A8989898989898888888888888787878787878686868686),
    .INIT_05(256'h909090908F8F8F8F8F8F8E8E8E8E8E8E8D8D8D8D8D8D8C8C8C8C8C8C8B8B8B8B),
    .INIT_06(256'h9595959595949494949494939393939393929292929292919191919191909090),
    .INIT_07(256'h9A9A9A9A9A9A9999999999999898989898989797979797979696969696969595),
    .INIT_08(256'h9F9F9F9F9F9F9E9E9E9E9E9E9E9D9D9D9D9D9D9C9C9C9C9C9C9B9B9B9B9B9B9A),
    .INIT_09(256'hA5A4A4A4A4A4A4A3A3A3A3A3A3A2A2A2A2A2A2A2A1A1A1A1A1A1A0A0A0A0A0A0),
    .INIT_0A(256'hAAAAA9A9A9A9A9A9A8A8A8A8A8A8A7A7A7A7A7A7A6A6A6A6A6A6A6A5A5A5A5A5),
    .INIT_0B(256'hAFAFAEAEAEAEAEAEADADADADADADADACACACACACACABABABABABABAAAAAAAAAA),
    .INIT_0C(256'hB4B4B4B3B3B3B3B3B3B2B2B2B2B2B2B1B1B1B1B1B1B1B0B0B0B0B0B0AFAFAFAF),
    .INIT_0D(256'hB9B9B9B8B8B8B8B8B8B7B7B7B7B7B7B7B6B6B6B6B6B6B5B5B5B5B5B5B4B4B4B4),
    .INIT_0E(256'hBEBEBEBEBDBDBDBDBDBDBCBCBCBCBCBCBBBBBBBBBBBBBBBABABABABABAB9B9B9),
    .INIT_0F(256'hC3C3C3C3C2C2C2C2C2C2C1C1C1C1C1C1C1C0C0C0C0C0C0BFBFBFBFBFBFBEBEBE),
    .INIT_10(256'hC8C8C8C8C7C7C7C7C7C7C7C6C6C6C6C6C6C5C5C5C5C5C5C4C4C4C4C4C4C4C3C3),
    .INIT_11(256'hCDCDCDCDCCCCCCCCCCCCCCCBCBCBCBCBCBCACACACACACAC9C9C9C9C9C9C9C8C8),
    .INIT_12(256'hD2D2D2D2D1D1D1D1D1D1D1D0D0D0D0D0D0CFCFCFCFCFCFCFCECECECECECECDCD),
    .INIT_13(256'hD7D7D7D7D7D6D6D6D6D6D6D5D5D5D5D5D5D4D4D4D4D4D4D4D3D3D3D3D3D3D2D2),
    .INIT_14(256'hDCDCDCDCDBDBDBDBDBDBDBDADADADADADAD9D9D9D9D9D9D9D8D8D8D8D8D8D7D7),
    .INIT_15(256'hE1E1E1E1E0E0E0E0E0E0E0DFDFDFDFDFDFDEDEDEDEDEDEDEDDDDDDDDDDDDDCDC),
    .INIT_16(256'hE6E6E6E6E5E5E5E5E5E5E5E4E4E4E4E4E4E3E3E3E3E3E3E3E2E2E2E2E2E2E1E1),
    .INIT_17(256'hEBEBEBEBEAEAEAEAEAEAE9E9E9E9E9E9E9E8E8E8E8E8E8E7E7E7E7E7E7E7E6E6),
    .INIT_18(256'hF0F0F0F0EFEFEFEFEFEFEEEEEEEEEEEEEEEDEDEDEDEDEDECECECECECECEBEBEB),
    .INIT_19(256'hF5F5F5F4F4F4F4F4F4F4F3F3F3F3F3F3F2F2F2F2F2F2F2F1F1F1F1F1F1F0F0F0),
    .INIT_1A(256'hFAFAFAF9F9F9F9F9F9F8F8F8F8F8F8F8F7F7F7F7F7F7F6F6F6F6F6F6F6F5F5F5),
    .INIT_1B(256'hFFFFFEFEFEFEFEFEFEFDFDFDFDFDFDFCFCFCFCFCFCFCFBFBFBFBFBFBFAFAFAFA),
    .INIT_1C(256'h04030303030303030202020202020201010101010100000000000000FFFFFFFF),
    .INIT_1D(256'h0908080808080807070707070707060606060606050505050505050404040404),
    .INIT_1E(256'h0D0D0D0D0D0D0C0C0C0C0C0C0C0B0B0B0B0B0B0B0A0A0A0A0A0A090909090909),
    .INIT_1F(256'h121212121212111111111111101010101010100F0F0F0F0F0F0E0E0E0E0E0E0E),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_055296_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_Naddra_o_al_n100 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i54_008,inst_doa_i54_007,inst_doa_i54_006,inst_doa_i54_005,inst_doa_i54_004,inst_doa_i54_003,inst_doa_i54_002,inst_doa_i54_001,inst_doa_i54_000}));
  // address_offset=56320;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'h1717171717161616161616151515151515151414141414141313131313131312),
    .INIT_01(256'h1C1C1C1C1B1B1B1B1B1B1A1A1A1A1A1A1A191919191919181818181818181717),
    .INIT_02(256'h2121202020202020201F1F1F1F1F1F1F1E1E1E1E1E1E1D1D1D1D1D1D1D1C1C1C),
    .INIT_03(256'h2625252525252525242424242424232323232323232222222222222221212121),
    .INIT_04(256'h2A2A2A2A2A2A2929292929292928282828282828272727272727262626262626),
    .INIT_05(256'h2F2F2F2F2F2E2E2E2E2E2E2E2D2D2D2D2D2D2C2C2C2C2C2C2C2B2B2B2B2B2B2B),
    .INIT_06(256'h3434343433333333333332323232323232313131313131313030303030302F2F),
    .INIT_07(256'h3939383838383838383737373737373636363636363635353535353535343434),
    .INIT_08(256'h3D3D3D3D3D3D3D3C3C3C3C3C3C3C3B3B3B3B3B3B3B3A3A3A3A3A3A3939393939),
    .INIT_09(256'h424242424241414141414141404040404040403F3F3F3F3F3F3F3E3E3E3E3E3E),
    .INIT_0A(256'h4747474646464646464645454545454545444444444444444343434343434342),
    .INIT_0B(256'h4C4C4B4B4B4B4B4B4A4A4A4A4A4A4A4949494949494948484848484848474747),
    .INIT_0C(256'h5050505050504F4F4F4F4F4F4F4E4E4E4E4E4E4E4D4D4D4D4D4D4D4C4C4C4C4C),
    .INIT_0D(256'h5555555554545454545454535353535353535252525252525251515151515150),
    .INIT_0E(256'h5A5A595959595959595858585858585857575757575756565656565656555555),
    .INIT_0F(256'h5E5E5E5E5E5E5D5D5D5D5D5D5D5C5C5C5C5C5C5C5B5B5B5B5B5B5B5A5A5A5A5A),
    .INIT_10(256'h636363636262626262626261616161616161606060606060605F5F5F5F5F5F5F),
    .INIT_11(256'h6868676767676767666666666666666565656565656564646464646464636363),
    .INIT_12(256'h6C6C6C6C6C6C6B6B6B6B6B6B6B6A6A6A6A6A6A6A696969696969696868686868),
    .INIT_13(256'h717171707070707070706F6F6F6F6F6F6F6E6E6E6E6E6E6E6D6D6D6D6D6D6D6C),
    .INIT_14(256'h7575757575757574747474747474737373737373737272727272727271717171),
    .INIT_15(256'h7A7A7A7A79797979797979787878787878787777777777777776767676767676),
    .INIT_16(256'h7F7E7E7E7E7E7E7E7D7D7D7D7D7D7D7C7C7C7C7C7C7C7B7B7B7B7B7B7B7A7A7A),
    .INIT_17(256'h83838383838282828282828281818181818181808080808080807F7F7F7F7F7F),
    .INIT_18(256'h8888878787878787878686868686868685858585858585848484848484848383),
    .INIT_19(256'h8C8C8C8C8C8C8B8B8B8B8B8B8B8A8A8A8A8A8A8A898989898989898888888888),
    .INIT_1A(256'h919191909090909090908F8F8F8F8F8F8F8E8E8E8E8E8E8E8D8D8D8D8D8D8D8C),
    .INIT_1B(256'h9595959595959494949494949493939393939393929292929292929191919191),
    .INIT_1C(256'h9A9A999999999999999998989898989898979797979797979696969696969695),
    .INIT_1D(256'h9E9E9E9E9E9E9D9D9D9D9D9D9D9C9C9C9C9C9C9C9B9B9B9B9B9B9B9A9A9A9A9A),
    .INIT_1E(256'hA3A3A2A2A2A2A2A2A2A1A1A1A1A1A1A1A0A0A0A0A0A0A0A09F9F9F9F9F9F9F9E),
    .INIT_1F(256'hA7A7A7A7A7A6A6A6A6A6A6A6A5A5A5A5A5A5A5A5A4A4A4A4A4A4A4A3A3A3A3A3),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_056320_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_Naddra_o_al_n100 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i55_008,inst_doa_i55_007,inst_doa_i55_006,inst_doa_i55_005,inst_doa_i55_004,inst_doa_i55_003,inst_doa_i55_002,inst_doa_i55_001,inst_doa_i55_000}));
  // address_offset=57344;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'h0000000000000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hACABABABABABABABAAAAAAAAAAAAAAAAA9A9A9A9A9A9A9A8A8A8A8A8A8A8A7A7),
    .INIT_01(256'hB0B0B0B0AFAFAFAFAFAFAFAFAEAEAEAEAEAEAEADADADADADADADACACACACACAC),
    .INIT_02(256'hB4B4B4B4B4B4B4B3B3B3B3B3B3B3B3B2B2B2B2B2B2B2B1B1B1B1B1B1B1B0B0B0),
    .INIT_03(256'hB9B9B9B8B8B8B8B8B8B8B7B7B7B7B7B7B7B6B6B6B6B6B6B6B6B5B5B5B5B5B5B5),
    .INIT_04(256'hBDBDBDBDBDBDBCBCBCBCBCBCBCBBBBBBBBBBBBBBBABABABABABABABAB9B9B9B9),
    .INIT_05(256'hC2C1C1C1C1C1C1C1C0C0C0C0C0C0C0C0BFBFBFBFBFBFBFBEBEBEBEBEBEBEBDBD),
    .INIT_06(256'hC6C6C6C6C5C5C5C5C5C5C5C4C4C4C4C4C4C4C3C3C3C3C3C3C3C3C2C2C2C2C2C2),
    .INIT_07(256'hCACACACACACAC9C9C9C9C9C9C9C8C8C8C8C8C8C8C8C7C7C7C7C7C7C7C6C6C6C6),
    .INIT_08(256'hCFCECECECECECECECECDCDCDCDCDCDCDCCCCCCCCCCCCCCCBCBCBCBCBCBCBCBCA),
    .INIT_09(256'hD3D3D3D2D2D2D2D2D2D2D2D1D1D1D1D1D1D1D0D0D0D0D0D0D0D0CFCFCFCFCFCF),
    .INIT_0A(256'hD7D7D7D7D7D7D6D6D6D6D6D6D6D5D5D5D5D5D5D5D5D4D4D4D4D4D4D4D3D3D3D3),
    .INIT_0B(256'hDBDBDBDBDBDBDBDBDADADADADADADAD9D9D9D9D9D9D9D9D8D8D8D8D8D8D8D7D7),
    .INIT_0C(256'hE0E0DFDFDFDFDFDFDFDFDEDEDEDEDEDEDEDDDDDDDDDDDDDDDDDCDCDCDCDCDCDC),
    .INIT_0D(256'hE4E4E4E4E3E3E3E3E3E3E3E3E2E2E2E2E2E2E2E1E1E1E1E1E1E1E1E0E0E0E0E0),
    .INIT_0E(256'hE8E8E8E8E8E8E7E7E7E7E7E7E7E7E6E6E6E6E6E6E6E5E5E5E5E5E5E5E5E4E4E4),
    .INIT_0F(256'hECECECECECECECECEBEBEBEBEBEBEBEAEAEAEAEAEAEAEAE9E9E9E9E9E9E9E9E8),
    .INIT_10(256'hF1F1F0F0F0F0F0F0F0EFEFEFEFEFEFEFEFEEEEEEEEEEEEEEEEEDEDEDEDEDEDED),
    .INIT_11(256'hF5F5F5F4F4F4F4F4F4F4F4F3F3F3F3F3F3F3F3F2F2F2F2F2F2F2F1F1F1F1F1F1),
    .INIT_12(256'hF9F9F9F9F9F8F8F8F8F8F8F8F7F7F7F7F7F7F7F7F6F6F6F6F6F6F6F6F5F5F5F5),
    .INIT_13(256'hFDFDFDFDFDFDFCFCFCFCFCFCFCFCFBFBFBFBFBFBFBFAFAFAFAFAFAFAFAF9F9F9),
    .INIT_14(256'h010101010101010000000000000000FFFFFFFFFFFFFFFFFEFEFEFEFEFEFEFDFD),
    .INIT_15(256'h0605050505050505040404040404040403030303030303030202020202020202),
    .INIT_16(256'h0A0A090909090909090808080808080808070707070707070706060606060606),
    .INIT_17(256'h0E0E0E0D0D0D0D0D0D0D0C0C0C0C0C0C0C0C0B0B0B0B0B0B0B0B0A0A0A0A0A0A),
    .INIT_18(256'h121212111111111111111110101010101010100F0F0F0F0F0F0F0F0E0E0E0E0E),
    .INIT_19(256'h1616161615151515151515151414141414141414131313131313131212121212),
    .INIT_1A(256'h1A1A1A1A19191919191919191818181818181818171717171717171716161616),
    .INIT_1B(256'h1E1E1E1E1E1D1D1D1D1D1D1D1D1C1C1C1C1C1C1C1C1B1B1B1B1B1B1B1B1A1A1A),
    .INIT_1C(256'h2222222222212121212121212120202020202020201F1F1F1F1F1F1F1F1E1E1E),
    .INIT_1D(256'h2626262626252525252525252524242424242424242323232323232323222222),
    .INIT_1E(256'h2A2A2A2A2A292929292929292928282828282828282727272727272727262626),
    .INIT_1F(256'h2E2E2E2E2E2D2D2D2D2D2D2D2D2C2C2C2C2C2C2C2C2B2B2B2B2B2B2B2B2A2A2A),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_057344_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_addra_o_al_n108 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i56_008,inst_doa_i56_007,inst_doa_i56_006,inst_doa_i56_005,inst_doa_i56_004,inst_doa_i56_003,inst_doa_i56_002,inst_doa_i56_001,inst_doa_i56_000}));
  // address_offset=57344;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000000000000000000000000000),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_057344_009 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n3504,open_n3505,open_n3506,open_n3507,open_n3508,open_n3509,open_n3510,1'b0,open_n3511}),
    .rsta(rsta),
    .doa({open_n3526,open_n3527,open_n3528,open_n3529,open_n3530,open_n3531,open_n3532,open_n3533,inst_doa_i56_009}));
  // address_offset=57344;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=12;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_057344_010 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa(addra[15:13]),
    .dia({open_n3562,open_n3563,open_n3564,open_n3565,open_n3566,open_n3567,open_n3568,1'b0,open_n3569}),
    .rsta(rsta),
    .doa({open_n3584,open_n3585,open_n3586,open_n3587,open_n3588,open_n3589,open_n3590,open_n3591,inst_doa_i56_010}));
  // address_offset=58368;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h3232323232313131313131313130303030303030302F2F2F2F2F2F2F2F2E2E2E),
    .INIT_01(256'h3636363636353535353535353534343434343434343333333333333333323232),
    .INIT_02(256'h3A3A3A3A3A393939393939393938383838383838383737373737373737363636),
    .INIT_03(256'h3E3E3E3E3D3D3D3D3D3D3D3D3C3C3C3C3C3C3C3C3B3B3B3B3B3B3B3B3A3A3A3A),
    .INIT_04(256'h42424241414141414141414140404040404040403F3F3F3F3F3F3F3F3E3E3E3E),
    .INIT_05(256'h4646464545454545454545444444444444444443434343434343434242424242),
    .INIT_06(256'h4A4A494949494949494948484848484848484747474747474747464646464646),
    .INIT_07(256'h4E4D4D4D4D4D4D4D4D4C4C4C4C4C4C4C4C4B4B4B4B4B4B4B4B4A4A4A4A4A4A4A),
    .INIT_08(256'h515151515151515150505050505050504F4F4F4F4F4F4F4F4E4E4E4E4E4E4E4E),
    .INIT_09(256'h5555555555555454545454545454545353535353535353525252525252525251),
    .INIT_0A(256'h5959595959585858585858585857575757575757575756565656565656565555),
    .INIT_0B(256'h5D5D5D5D5C5C5C5C5C5C5C5C5B5B5B5B5B5B5B5B5A5A5A5A5A5A5A5A5A595959),
    .INIT_0C(256'h616160606060606060605F5F5F5F5F5F5F5F5F5E5E5E5E5E5E5E5E5D5D5D5D5D),
    .INIT_0D(256'h6464646464646464636363636363636363626262626262626261616161616161),
    .INIT_0E(256'h6868686868686767676767676767676666666666666666656565656565656565),
    .INIT_0F(256'h6C6C6C6C6B6B6B6B6B6B6B6B6B6A6A6A6A6A6A6A6A6969696969696969696868),
    .INIT_10(256'h70706F6F6F6F6F6F6F6F6F6E6E6E6E6E6E6E6E6D6D6D6D6D6D6D6D6D6C6C6C6C),
    .INIT_11(256'h7373737373737373727272727272727272717171717171717171707070707070),
    .INIT_12(256'h7777777777777676767676767676757575757575757575747474747474747474),
    .INIT_13(256'h7B7B7B7A7A7A7A7A7A7A7A7A7979797979797979787878787878787878777777),
    .INIT_14(256'h7E7E7E7E7E7E7E7E7E7D7D7D7D7D7D7D7D7D7C7C7C7C7C7C7C7C7B7B7B7B7B7B),
    .INIT_15(256'h82828282828281818181818181818180808080808080807F7F7F7F7F7F7F7F7F),
    .INIT_16(256'h8686868585858585858585858484848484848484838383838383838383828282),
    .INIT_17(256'h8989898989898989888888888888888888878787878787878787868686868686),
    .INIT_18(256'h8D8D8D8D8D8C8C8C8C8C8C8C8C8C8B8B8B8B8B8B8B8B8B8A8A8A8A8A8A8A8A8A),
    .INIT_19(256'h919090909090909090908F8F8F8F8F8F8F8F8F8E8E8E8E8E8E8E8E8E8D8D8D8D),
    .INIT_1A(256'h9494949494949493939393939393939292929292929292929191919191919191),
    .INIT_1B(256'h9898989797979797979797979696969696969696969595959595959595959494),
    .INIT_1C(256'h9B9B9B9B9B9B9B9B9A9A9A9A9A9A9A9A9A999999999999999999989898989898),
    .INIT_1D(256'h9F9F9F9E9E9E9E9E9E9E9E9E9D9D9D9D9D9D9D9D9D9C9C9C9C9C9C9C9C9C9C9B),
    .INIT_1E(256'hA2A2A2A2A2A2A2A2A1A1A1A1A1A1A1A1A1A0A0A0A0A0A0A0A0A09F9F9F9F9F9F),
    .INIT_1F(256'hA6A6A6A5A5A5A5A5A5A5A5A5A5A4A4A4A4A4A4A4A4A4A3A3A3A3A3A3A3A3A3A2),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_058368_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_addra_o_al_n108 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i57_008,inst_doa_i57_007,inst_doa_i57_006,inst_doa_i57_005,inst_doa_i57_004,inst_doa_i57_003,inst_doa_i57_002,inst_doa_i57_001,inst_doa_i57_000}));
  // address_offset=59392;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000000000000000000000),
    .INIT_00(256'hA9A9A9A9A9A9A9A9A8A8A8A8A8A8A8A8A8A7A7A7A7A7A7A7A7A7A6A6A6A6A6A6),
    .INIT_01(256'hADADADACACACACACACACACACABABABABABABABABABABAAAAAAAAAAAAAAAAAAA9),
    .INIT_02(256'hB0B0B0B0B0B0B0AFAFAFAFAFAFAFAFAFAFAEAEAEAEAEAEAEAEAEADADADADADAD),
    .INIT_03(256'hB4B4B3B3B3B3B3B3B3B3B3B2B2B2B2B2B2B2B2B2B2B1B1B1B1B1B1B1B1B1B0B0),
    .INIT_04(256'hB7B7B7B7B7B7B6B6B6B6B6B6B6B6B6B5B5B5B5B5B5B5B5B5B5B4B4B4B4B4B4B4),
    .INIT_05(256'hBABABABABABABABABABAB9B9B9B9B9B9B9B9B9B8B8B8B8B8B8B8B8B8B8B7B7B7),
    .INIT_06(256'hBEBEBEBEBDBDBDBDBDBDBDBDBDBCBCBCBCBCBCBCBCBCBCBBBBBBBBBBBBBBBBBB),
    .INIT_07(256'hC1C1C1C1C1C1C1C0C0C0C0C0C0C0C0C0C0BFBFBFBFBFBFBFBFBFBEBEBEBEBEBE),
    .INIT_08(256'hC5C4C4C4C4C4C4C4C4C4C4C3C3C3C3C3C3C3C3C3C2C2C2C2C2C2C2C2C2C2C1C1),
    .INIT_09(256'hC8C8C8C8C8C7C7C7C7C7C7C7C7C7C6C6C6C6C6C6C6C6C6C6C5C5C5C5C5C5C5C5),
    .INIT_0A(256'hCBCBCBCBCBCBCBCBCACACACACACACACACAC9C9C9C9C9C9C9C9C9C9C8C8C8C8C8),
    .INIT_0B(256'hCFCECECECECECECECECECECDCDCDCDCDCDCDCDCDCCCCCCCCCCCCCCCCCCCCCBCB),
    .INIT_0C(256'hD2D2D2D2D1D1D1D1D1D1D1D1D1D1D0D0D0D0D0D0D0D0D0CFCFCFCFCFCFCFCFCF),
    .INIT_0D(256'hD5D5D5D5D5D5D4D4D4D4D4D4D4D4D4D4D3D3D3D3D3D3D3D3D3D3D2D2D2D2D2D2),
    .INIT_0E(256'hD8D8D8D8D8D8D8D8D8D7D7D7D7D7D7D7D7D7D7D6D6D6D6D6D6D6D6D6D6D5D5D5),
    .INIT_0F(256'hDCDBDBDBDBDBDBDBDBDBDBDADADADADADADADADADAD9D9D9D9D9D9D9D9D9D9D8),
    .INIT_10(256'hDFDFDFDFDEDEDEDEDEDEDEDEDEDEDDDDDDDDDDDDDDDDDDDDDCDCDCDCDCDCDCDC),
    .INIT_11(256'hE2E2E2E2E2E2E1E1E1E1E1E1E1E1E1E1E0E0E0E0E0E0E0E0E0E0DFDFDFDFDFDF),
    .INIT_12(256'hE5E5E5E5E5E5E5E5E4E4E4E4E4E4E4E4E4E4E3E3E3E3E3E3E3E3E3E3E2E2E2E2),
    .INIT_13(256'hE8E8E8E8E8E8E8E8E8E7E7E7E7E7E7E7E7E7E7E7E6E6E6E6E6E6E6E6E6E6E5E5),
    .INIT_14(256'hECEBEBEBEBEBEBEBEBEBEBEAEAEAEAEAEAEAEAEAEAE9E9E9E9E9E9E9E9E9E9E8),
    .INIT_15(256'hEFEFEEEEEEEEEEEEEEEEEEEEEEEDEDEDEDEDEDEDEDEDEDECECECECECECECECEC),
    .INIT_16(256'hF2F2F2F2F1F1F1F1F1F1F1F1F1F1F0F0F0F0F0F0F0F0F0F0EFEFEFEFEFEFEFEF),
    .INIT_17(256'hF5F5F5F5F5F4F4F4F4F4F4F4F4F4F4F3F3F3F3F3F3F3F3F3F3F2F2F2F2F2F2F2),
    .INIT_18(256'hF8F8F8F8F8F8F7F7F7F7F7F7F7F7F7F7F6F6F6F6F6F6F6F6F6F6F5F5F5F5F5F5),
    .INIT_19(256'hFBFBFBFBFBFBFAFAFAFAFAFAFAFAFAFAFAF9F9F9F9F9F9F9F9F9F9F8F8F8F8F8),
    .INIT_1A(256'hFEFEFEFEFEFEFEFDFDFDFDFDFDFDFDFDFDFDFCFCFCFCFCFCFCFCFCFCFBFBFBFB),
    .INIT_1B(256'h010101010101010000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFEFEFE),
    .INIT_1C(256'h0404040404040404030303030303030303030202020202020202020202010101),
    .INIT_1D(256'h0707070707070707060606060606060606060505050505050505050505040404),
    .INIT_1E(256'h0A0A0A0A0A0A0A0A090909090909090909090808080808080808080808070707),
    .INIT_1F(256'h0D0D0D0D0D0D0D0C0C0C0C0C0C0C0C0C0C0C0B0B0B0B0B0B0B0B0B0B0B0A0A0A),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_059392_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_addra_o_al_n108 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i58_008,inst_doa_i58_007,inst_doa_i58_006,inst_doa_i58_005,inst_doa_i58_004,inst_doa_i58_003,inst_doa_i58_002,inst_doa_i58_001,inst_doa_i58_000}));
  // address_offset=60416;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'h101010101010100F0F0F0F0F0F0F0F0F0F0F0E0E0E0E0E0E0E0E0E0E0E0D0D0D),
    .INIT_01(256'h1313131313131212121212121212121212111111111111111111111110101010),
    .INIT_02(256'h1616161616151515151515151515151514141414141414141414141313131313),
    .INIT_03(256'h1919191918181818181818181818181717171717171717171717161616161616),
    .INIT_04(256'h1C1C1C1B1B1B1B1B1B1B1B1B1B1B1A1A1A1A1A1A1A1A1A1A1A19191919191919),
    .INIT_05(256'h1F1F1E1E1E1E1E1E1E1E1E1E1E1D1D1D1D1D1D1D1D1D1D1D1C1C1C1C1C1C1C1C),
    .INIT_06(256'h212121212121212121212120202020202020202020201F1F1F1F1F1F1F1F1F1F),
    .INIT_07(256'h2424242424242424242323232323232323232323232222222222222222222222),
    .INIT_08(256'h2727272727272726262626262626262626262625252525252525252525252424),
    .INIT_09(256'h2A2A2A2A2A292929292929292929292929282828282828282828282827272727),
    .INIT_0A(256'h2D2D2D2C2C2C2C2C2C2C2C2C2C2C2B2B2B2B2B2B2B2B2B2B2B2B2A2A2A2A2A2A),
    .INIT_0B(256'h2F2F2F2F2F2F2F2F2F2F2F2F2E2E2E2E2E2E2E2E2E2E2E2D2D2D2D2D2D2D2D2D),
    .INIT_0C(256'h3232323232323232323131313131313131313131303030303030303030303030),
    .INIT_0D(256'h3535353535353434343434343434343434333333333333333333333333323232),
    .INIT_0E(256'h3838373737373737373737373737363636363636363636363636353535353535),
    .INIT_0F(256'h3A3A3A3A3A3A3A3A3A3A39393939393939393939393938383838383838383838),
    .INIT_10(256'h3D3D3D3D3D3D3D3C3C3C3C3C3C3C3C3C3C3C3C3B3B3B3B3B3B3B3B3B3B3B3B3A),
    .INIT_11(256'h4040403F3F3F3F3F3F3F3F3F3F3F3F3E3E3E3E3E3E3E3E3E3E3E3E3D3D3D3D3D),
    .INIT_12(256'h4242424242424242424241414141414141414141414140404040404040404040),
    .INIT_13(256'h4545454545454444444444444444444444444343434343434343434343434242),
    .INIT_14(256'h4847474747474747474747474746464646464646464646464646454545454545),
    .INIT_15(256'h4A4A4A4A4A4A4A4A494949494949494949494949494848484848484848484848),
    .INIT_16(256'h4D4D4D4C4C4C4C4C4C4C4C4C4C4C4C4C4B4B4B4B4B4B4B4B4B4B4B4B4A4A4A4A),
    .INIT_17(256'h4F4F4F4F4F4F4F4F4F4F4E4E4E4E4E4E4E4E4E4E4E4E4E4D4D4D4D4D4D4D4D4D),
    .INIT_18(256'h5252525251515151515151515151515151505050505050505050505050504F4F),
    .INIT_19(256'h5454545454545454545454535353535353535353535353535252525252525252),
    .INIT_1A(256'h5757575757565656565656565656565656555555555555555555555555555454),
    .INIT_1B(256'h5959595959595959595959585858585858585858585858585757575757575757),
    .INIT_1C(256'h5C5C5C5C5B5B5B5B5B5B5B5B5B5B5B5B5B5A5A5A5A5A5A5A5A5A5A5A5A5A5959),
    .INIT_1D(256'h5E5E5E5E5E5E5E5E5E5E5D5D5D5D5D5D5D5D5D5D5D5D5D5C5C5C5C5C5C5C5C5C),
    .INIT_1E(256'h616161606060606060606060606060605F5F5F5F5F5F5F5F5F5F5F5F5F5E5E5E),
    .INIT_1F(256'h6363636363636363626262626262626262626262626161616161616161616161),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_060416_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_Naddra[12]_addra_o_al_n108 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i59_008,inst_doa_i59_007,inst_doa_i59_006,inst_doa_i59_005,inst_doa_i59_004,inst_doa_i59_003,inst_doa_i59_002,inst_doa_i59_001,inst_doa_i59_000}));
  // address_offset=61440;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'h6565656565656565656565656564646464646464646464646464646363636363),
    .INIT_01(256'h6868686868676767676767676767676767676766666666666666666666666666),
    .INIT_02(256'h6A6A6A6A6A6A6A6A6A6A69696969696969696969696969696868686868686868),
    .INIT_03(256'h6D6C6C6C6C6C6C6C6C6C6C6C6C6C6C6B6B6B6B6B6B6B6B6B6B6B6B6B6A6A6A6A),
    .INIT_04(256'h6F6F6F6F6F6F6E6E6E6E6E6E6E6E6E6E6E6E6E6D6D6D6D6D6D6D6D6D6D6D6D6D),
    .INIT_05(256'h7171717171717171717170707070707070707070707070706F6F6F6F6F6F6F6F),
    .INIT_06(256'h7373737373737373737373737373727272727272727272727272727271717171),
    .INIT_07(256'h7676767675757575757575757575757575757474747474747474747474747474),
    .INIT_08(256'h7878787878787877777777777777777777777777777776767676767676767676),
    .INIT_09(256'h7A7A7A7A7A7A7A7A7A7A7A797979797979797979797979797978787878787878),
    .INIT_0A(256'h7C7C7C7C7C7C7C7C7C7C7C7C7C7C7B7B7B7B7B7B7B7B7B7B7B7B7B7B7A7A7A7A),
    .INIT_0B(256'h7F7F7E7E7E7E7E7E7E7E7E7E7E7E7E7E7E7D7D7D7D7D7D7D7D7D7D7D7D7D7D7D),
    .INIT_0C(256'h81818181818080808080808080808080808080807F7F7F7F7F7F7F7F7F7F7F7F),
    .INIT_0D(256'h8383838383838383828282828282828282828282828281818181818181818181),
    .INIT_0E(256'h8585858585858585858584848484848484848484848484848483838383838383),
    .INIT_0F(256'h8787878787878787878787878686868686868686868686868686868585858585),
    .INIT_10(256'h8989898989898989898989898988888888888888888888888888888888878787),
    .INIT_11(256'h8B8B8B8B8B8B8B8B8B8B8B8B8B8B8B8A8A8A8A8A8A8A8A8A8A8A8A8A8A8A8989),
    .INIT_12(256'h8E8D8D8D8D8D8D8D8D8D8D8D8D8D8D8D8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C),
    .INIT_13(256'h90908F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8E8E8E8E8E8E8E8E8E8E8E8E8E8E8E),
    .INIT_14(256'h9292919191919191919191919191919191919090909090909090909090909090),
    .INIT_15(256'h9494939393939393939393939393939393939292929292929292929292929292),
    .INIT_16(256'h9696959595959595959595959595959595959494949494949494949494949494),
    .INIT_17(256'h9898979797979797979797979797979797979696969696969696969696969696),
    .INIT_18(256'h9A99999999999999999999999999999999999898989898989898989898989898),
    .INIT_19(256'h9C9B9B9B9B9B9B9B9B9B9B9B9B9B9B9B9B9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A),
    .INIT_1A(256'h9D9D9D9D9D9D9D9D9D9D9D9D9D9D9D9D9C9C9C9C9C9C9C9C9C9C9C9C9C9C9C9C),
    .INIT_1B(256'h9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9E9E9E9E9E9E9E9E9E9E9E9E9E9E9E9E9D),
    .INIT_1C(256'hA1A1A1A1A1A1A1A1A1A1A1A1A1A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A09F9F),
    .INIT_1D(256'hA3A3A3A3A3A3A3A3A3A3A3A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A2A1A1A1A1),
    .INIT_1E(256'hA5A5A5A5A5A5A5A5A4A4A4A4A4A4A4A4A4A4A4A4A4A4A4A4A4A4A3A3A3A3A3A3),
    .INIT_1F(256'hA7A7A7A7A7A6A6A6A6A6A6A6A6A6A6A6A6A6A6A6A6A6A6A5A5A5A5A5A5A5A5A5),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_061440_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_addra[_o_al_n116 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i60_008,inst_doa_i60_007,inst_doa_i60_006,inst_doa_i60_005,inst_doa_i60_004,inst_doa_i60_003,inst_doa_i60_002,inst_doa_i60_001,inst_doa_i60_000}));
  // address_offset=62464;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'hA9A9A8A8A8A8A8A8A8A8A8A8A8A8A8A8A8A8A8A8A7A7A7A7A7A7A7A7A7A7A7A7),
    .INIT_01(256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9A9A9A9A9A9A9A9A9A9A9A9A9A9A9A9),
    .INIT_02(256'hACACACACACACACACACACACACACABABABABABABABABABABABABABABABABABABAA),
    .INIT_03(256'hAEAEAEAEAEAEAEAEADADADADADADADADADADADADADADADADADADACACACACACAC),
    .INIT_04(256'hB0B0B0B0AFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAEAEAEAEAEAEAEAEAEAE),
    .INIT_05(256'hB1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B1B0B0B0B0B0B0B0B0B0B0B0B0B0B0B0),
    .INIT_06(256'hB3B3B3B3B3B3B3B3B3B3B3B3B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B2B1B1),
    .INIT_07(256'hB5B5B5B5B5B5B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B4B3B3B3B3B3B3B3),
    .INIT_08(256'hB6B6B6B6B6B6B6B6B6B6B6B6B6B6B6B6B6B6B6B5B5B5B5B5B5B5B5B5B5B5B5B5),
    .INIT_09(256'hB8B8B8B8B8B8B8B8B8B8B8B8B7B7B7B7B7B7B7B7B7B7B7B7B7B7B7B7B7B7B7B6),
    .INIT_0A(256'hBABABABABAB9B9B9B9B9B9B9B9B9B9B9B9B9B9B9B9B9B9B9B9B8B8B8B8B8B8B8),
    .INIT_0B(256'hBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBABABABABABABABABABABABABABABA),
    .INIT_0C(256'hBDBDBDBDBDBDBDBDBDBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBBBBBB),
    .INIT_0D(256'hBFBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBDBDBDBDBDBDBDBDBDBDBD),
    .INIT_0E(256'hC0C0C0C0C0C0C0C0C0C0C0C0BFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBF),
    .INIT_0F(256'hC2C2C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C1C0C0C0C0C0C0C0C0C0),
    .INIT_10(256'hC3C3C3C3C3C3C3C3C3C3C3C3C3C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2C2),
    .INIT_11(256'hC5C5C5C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C4C3C3C3C3C3C3C3C3),
    .INIT_12(256'hC6C6C6C6C6C6C6C6C6C6C6C6C6C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5C5),
    .INIT_13(256'hC8C8C7C7C7C7C7C7C7C7C7C7C7C7C7C7C7C7C7C7C7C7C7C7C6C6C6C6C6C6C6C6),
    .INIT_14(256'hC9C9C9C9C9C9C9C9C9C9C9C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8C8),
    .INIT_15(256'hCACACACACACACACACACACACACACACACACACACACACAC9C9C9C9C9C9C9C9C9C9C9),
    .INIT_16(256'hCCCCCCCCCCCCCCCCCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCBCA),
    .INIT_17(256'hCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCCCCCCCCCCCCCCCCCCCCCCCCCCCCCC),
    .INIT_18(256'hCFCFCECECECECECECECECECECECECECECECECECECECECECECECECDCDCDCDCDCD),
    .INIT_19(256'hD0D0D0D0D0D0D0D0D0D0D0CFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCF),
    .INIT_1A(256'hD1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D1D0D0D0D0D0D0D0D0D0D0D0D0D0),
    .INIT_1B(256'hD3D3D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D2D1D1D1D1D1),
    .INIT_1C(256'hD4D4D4D4D4D4D4D4D4D3D3D3D3D3D3D3D3D3D3D3D3D3D3D3D3D3D3D3D3D3D3D3),
    .INIT_1D(256'hD5D5D5D5D5D5D5D5D5D5D5D5D5D5D5D5D4D4D4D4D4D4D4D4D4D4D4D4D4D4D4D4),
    .INIT_1E(256'hD6D6D6D6D6D6D6D6D6D6D6D6D6D6D6D6D6D6D6D6D6D6D6D5D5D5D5D5D5D5D5D5),
    .INIT_1F(256'hD8D8D8D8D7D7D7D7D7D7D7D7D7D7D7D7D7D7D7D7D7D7D7D7D7D7D7D7D7D7D6D6),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_062464_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_addra[_o_al_n116 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i61_008,inst_doa_i61_007,inst_doa_i61_006,inst_doa_i61_005,inst_doa_i61_004,inst_doa_i61_003,inst_doa_i61_002,inst_doa_i61_001,inst_doa_i61_000}));
  // address_offset=63488;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'hD9D9D9D9D9D9D9D9D9D8D8D8D8D8D8D8D8D8D8D8D8D8D8D8D8D8D8D8D8D8D8D8),
    .INIT_01(256'hDADADADADADADADADADADADADADADAD9D9D9D9D9D9D9D9D9D9D9D9D9D9D9D9D9),
    .INIT_02(256'hDBDBDBDBDBDBDBDBDBDBDBDBDBDBDBDBDBDBDBDBDADADADADADADADADADADADA),
    .INIT_03(256'hDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDCDBDBDBDBDBDBDB),
    .INIT_04(256'hDEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDCDCDC),
    .INIT_05(256'hDFDFDFDFDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDE),
    .INIT_06(256'hE0E0E0E0E0E0E0DFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDF),
    .INIT_07(256'hE1E1E1E1E1E1E1E1E1E1E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0E0),
    .INIT_08(256'hE2E2E2E2E2E2E2E2E2E2E2E2E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1E1),
    .INIT_09(256'hE3E3E3E3E3E3E3E3E3E3E3E3E3E3E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2E2),
    .INIT_0A(256'hE4E4E4E4E4E4E4E4E4E4E4E4E4E4E4E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3E3),
    .INIT_0B(256'hE5E5E5E5E5E5E5E5E5E5E5E5E5E5E5E4E4E4E4E4E4E4E4E4E4E4E4E4E4E4E4E4),
    .INIT_0C(256'hE6E6E6E6E6E6E6E6E6E6E6E6E6E6E6E5E5E5E5E5E5E5E5E5E5E5E5E5E5E5E5E5),
    .INIT_0D(256'hE7E7E7E7E7E7E7E7E7E7E7E7E7E7E7E6E6E6E6E6E6E6E6E6E6E6E6E6E6E6E6E6),
    .INIT_0E(256'hE8E8E8E8E8E8E8E8E8E8E8E8E8E7E7E7E7E7E7E7E7E7E7E7E7E7E7E7E7E7E7E7),
    .INIT_0F(256'hE9E9E9E9E9E9E9E9E9E9E9E8E8E8E8E8E8E8E8E8E8E8E8E8E8E8E8E8E8E8E8E8),
    .INIT_10(256'hEAEAEAEAEAEAEAEAE9E9E9E9E9E9E9E9E9E9E9E9E9E9E9E9E9E9E9E9E9E9E9E9),
    .INIT_11(256'hEBEBEBEBEBEAEAEAEAEAEAEAEAEAEAEAEAEAEAEAEAEAEAEAEAEAEAEAEAEAEAEA),
    .INIT_12(256'hEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEBEB),
    .INIT_13(256'hECECECECECECECECECECECECECECECECECECECECECECECECECECECECECECECEC),
    .INIT_14(256'hEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDEDECECECECEC),
    .INIT_15(256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEDEDEDEDEDEDEDEDEDEDEDED),
    .INIT_16(256'hEFEFEFEFEFEFEFEFEFEFEFEFEFEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE),
    .INIT_17(256'hF0F0F0F0EFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEF),
    .INIT_18(256'hF0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0),
    .INIT_19(256'hF1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F0F0F0F0F0F0),
    .INIT_1A(256'hF2F2F2F2F2F2F2F2F2F2F2F2F2F2F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1F1),
    .INIT_1B(256'hF3F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2F2),
    .INIT_1C(256'hF3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3F3),
    .INIT_1D(256'hF4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F3F3F3F3F3F3F3F3F3F3F3F3F3F3),
    .INIT_1E(256'hF4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4F4),
    .INIT_1F(256'hF5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_063488_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_addra[_o_al_n116 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i62_008,inst_doa_i62_007,inst_doa_i62_006,inst_doa_i62_005,inst_doa_i62_004,inst_doa_i62_003,inst_doa_i62_002,inst_doa_i62_001,inst_doa_i62_000}));
  // address_offset=64512;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=12;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INITP_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_00(256'hF6F6F6F6F6F6F6F6F6F6F6F6F6F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5F5),
    .INIT_01(256'hF6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6F6),
    .INIT_02(256'hF7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F6F6F6F6F6F6F6F6F6F6),
    .INIT_03(256'hF7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7F7),
    .INIT_04(256'hF8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F7F7F7),
    .INIT_05(256'hF8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8),
    .INIT_06(256'hF9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F8),
    .INIT_07(256'hF9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9F9),
    .INIT_08(256'hFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAF9F9F9F9),
    .INIT_09(256'hFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFAFA),
    .INIT_0A(256'hFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFAFAFAFAFAFAFAFAFAFAFAFAFA),
    .INIT_0B(256'hFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFB),
    .INIT_0C(256'hFCFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFBFB),
    .INIT_0D(256'hFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFC),
    .INIT_0E(256'hFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFC),
    .INIT_0F(256'hFDFDFDFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFCFC),
    .INIT_10(256'hFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFD),
    .INIT_11(256'hFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFD),
    .INIT_12(256'hFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFD),
    .INIT_13(256'hFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFDFD),
    .INIT_14(256'hFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE),
    .INIT_15(256'hFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE),
    .INIT_16(256'hFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE),
    .INIT_17(256'hFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE),
    .INIT_18(256'hFFFFFFFFFFFFFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFE),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_65536x12_sub_064512_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa({\and_addra[12]_addra[_o_al_n116 ,addra[11:10]}),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i63_008,inst_doa_i63_007,inst_doa_i63_006,inst_doa_i63_005,inst_doa_i63_004,inst_doa_i63_003,inst_doa_i63_002,inst_doa_i63_001,inst_doa_i63_000}));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_0  (
    .i0(inst_doa_i0_000),
    .i1(inst_doa_i1_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_0 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_1  (
    .i0(inst_doa_i2_000),
    .i1(inst_doa_i3_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_1 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_10  (
    .i0(inst_doa_i20_000),
    .i1(inst_doa_i21_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_10 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_11  (
    .i0(inst_doa_i22_000),
    .i1(inst_doa_i23_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_11 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_12  (
    .i0(inst_doa_i24_000),
    .i1(inst_doa_i25_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_12 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_13  (
    .i0(inst_doa_i26_000),
    .i1(inst_doa_i27_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_13 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_14  (
    .i0(inst_doa_i28_000),
    .i1(inst_doa_i29_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_14 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_15  (
    .i0(inst_doa_i30_000),
    .i1(inst_doa_i31_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_15 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_16  (
    .i0(inst_doa_i32_000),
    .i1(inst_doa_i33_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_16 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_17  (
    .i0(inst_doa_i34_000),
    .i1(inst_doa_i35_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_17 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_18  (
    .i0(inst_doa_i36_000),
    .i1(inst_doa_i37_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_18 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_19  (
    .i0(inst_doa_i38_000),
    .i1(inst_doa_i39_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_19 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_2  (
    .i0(inst_doa_i4_000),
    .i1(inst_doa_i5_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_2 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_20  (
    .i0(inst_doa_i40_000),
    .i1(inst_doa_i41_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_20 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_21  (
    .i0(inst_doa_i42_000),
    .i1(inst_doa_i43_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_21 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_22  (
    .i0(inst_doa_i44_000),
    .i1(inst_doa_i45_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_22 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_23  (
    .i0(inst_doa_i46_000),
    .i1(inst_doa_i47_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_23 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_24  (
    .i0(inst_doa_i48_000),
    .i1(inst_doa_i49_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_24 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_25  (
    .i0(inst_doa_i50_000),
    .i1(inst_doa_i51_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_25 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_26  (
    .i0(inst_doa_i52_000),
    .i1(inst_doa_i53_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_26 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_27  (
    .i0(inst_doa_i54_000),
    .i1(inst_doa_i55_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_27 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_28  (
    .i0(inst_doa_i56_000),
    .i1(inst_doa_i57_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_28 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_29  (
    .i0(inst_doa_i58_000),
    .i1(inst_doa_i59_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_29 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_3  (
    .i0(inst_doa_i6_000),
    .i1(inst_doa_i7_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_3 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_30  (
    .i0(inst_doa_i60_000),
    .i1(inst_doa_i61_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_30 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_31  (
    .i0(inst_doa_i62_000),
    .i1(inst_doa_i63_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_31 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_4  (
    .i0(inst_doa_i8_000),
    .i1(inst_doa_i9_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_4 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_5  (
    .i0(inst_doa_i10_000),
    .i1(inst_doa_i11_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_5 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_6  (
    .i0(inst_doa_i12_000),
    .i1(inst_doa_i13_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_6 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_7  (
    .i0(inst_doa_i14_000),
    .i1(inst_doa_i15_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_7 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_8  (
    .i0(inst_doa_i16_000),
    .i1(inst_doa_i17_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_8 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_9  (
    .i0(inst_doa_i18_000),
    .i1(inst_doa_i19_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_9 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b0/B0_0 ),
    .i1(\inst_doa_mux_b0/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_0 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b0/B0_2 ),
    .i1(\inst_doa_mux_b0/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_1 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_10  (
    .i0(\inst_doa_mux_b0/B0_20 ),
    .i1(\inst_doa_mux_b0/B0_21 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_10 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_11  (
    .i0(\inst_doa_mux_b0/B0_22 ),
    .i1(\inst_doa_mux_b0/B0_23 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_11 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_12  (
    .i0(\inst_doa_mux_b0/B0_24 ),
    .i1(\inst_doa_mux_b0/B0_25 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_12 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_13  (
    .i0(\inst_doa_mux_b0/B0_26 ),
    .i1(\inst_doa_mux_b0/B0_27 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_13 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_14  (
    .i0(\inst_doa_mux_b0/B0_28 ),
    .i1(\inst_doa_mux_b0/B0_29 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_14 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_15  (
    .i0(\inst_doa_mux_b0/B0_30 ),
    .i1(\inst_doa_mux_b0/B0_31 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_15 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_2  (
    .i0(\inst_doa_mux_b0/B0_4 ),
    .i1(\inst_doa_mux_b0/B0_5 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_2 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_3  (
    .i0(\inst_doa_mux_b0/B0_6 ),
    .i1(\inst_doa_mux_b0/B0_7 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_3 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_4  (
    .i0(\inst_doa_mux_b0/B0_8 ),
    .i1(\inst_doa_mux_b0/B0_9 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_4 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_5  (
    .i0(\inst_doa_mux_b0/B0_10 ),
    .i1(\inst_doa_mux_b0/B0_11 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_5 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_6  (
    .i0(\inst_doa_mux_b0/B0_12 ),
    .i1(\inst_doa_mux_b0/B0_13 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_6 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_7  (
    .i0(\inst_doa_mux_b0/B0_14 ),
    .i1(\inst_doa_mux_b0/B0_15 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_7 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_8  (
    .i0(\inst_doa_mux_b0/B0_16 ),
    .i1(\inst_doa_mux_b0/B0_17 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_8 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_9  (
    .i0(\inst_doa_mux_b0/B0_18 ),
    .i1(\inst_doa_mux_b0/B0_19 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_9 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b0/B1_0 ),
    .i1(\inst_doa_mux_b0/B1_1 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b0/B2_0 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_2_1  (
    .i0(\inst_doa_mux_b0/B1_2 ),
    .i1(\inst_doa_mux_b0/B1_3 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b0/B2_1 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_2_2  (
    .i0(\inst_doa_mux_b0/B1_4 ),
    .i1(\inst_doa_mux_b0/B1_5 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b0/B2_2 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_2_3  (
    .i0(\inst_doa_mux_b0/B1_6 ),
    .i1(\inst_doa_mux_b0/B1_7 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b0/B2_3 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_2_4  (
    .i0(\inst_doa_mux_b0/B1_8 ),
    .i1(\inst_doa_mux_b0/B1_9 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b0/B2_4 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_2_5  (
    .i0(\inst_doa_mux_b0/B1_10 ),
    .i1(\inst_doa_mux_b0/B1_11 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b0/B2_5 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_2_6  (
    .i0(\inst_doa_mux_b0/B1_12 ),
    .i1(\inst_doa_mux_b0/B1_13 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b0/B2_6 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_2_7  (
    .i0(\inst_doa_mux_b0/B1_14 ),
    .i1(\inst_doa_mux_b0/B1_15 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b0/B2_7 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_3_0  (
    .i0(\inst_doa_mux_b0/B2_0 ),
    .i1(\inst_doa_mux_b0/B2_1 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b0/B3_0 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_3_1  (
    .i0(\inst_doa_mux_b0/B2_2 ),
    .i1(\inst_doa_mux_b0/B2_3 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b0/B3_1 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_3_2  (
    .i0(\inst_doa_mux_b0/B2_4 ),
    .i1(\inst_doa_mux_b0/B2_5 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b0/B3_2 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_3_3  (
    .i0(\inst_doa_mux_b0/B2_6 ),
    .i1(\inst_doa_mux_b0/B2_7 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b0/B3_3 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_4_0  (
    .i0(\inst_doa_mux_b0/B3_0 ),
    .i1(\inst_doa_mux_b0/B3_1 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b0/B4_0 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_4_1  (
    .i0(\inst_doa_mux_b0/B3_2 ),
    .i1(\inst_doa_mux_b0/B3_3 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b0/B4_1 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_5_0  (
    .i0(\inst_doa_mux_b0/B4_0 ),
    .i1(\inst_doa_mux_b0/B4_1 ),
    .sel(addra_piped[5]),
    .o(doa[0]));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_0  (
    .i0(inst_doa_i0_001),
    .i1(inst_doa_i1_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_0 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_1  (
    .i0(inst_doa_i2_001),
    .i1(inst_doa_i3_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_1 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_10  (
    .i0(inst_doa_i20_001),
    .i1(inst_doa_i21_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_10 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_11  (
    .i0(inst_doa_i22_001),
    .i1(inst_doa_i23_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_11 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_12  (
    .i0(inst_doa_i24_001),
    .i1(inst_doa_i25_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_12 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_13  (
    .i0(inst_doa_i26_001),
    .i1(inst_doa_i27_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_13 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_14  (
    .i0(inst_doa_i28_001),
    .i1(inst_doa_i29_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_14 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_15  (
    .i0(inst_doa_i30_001),
    .i1(inst_doa_i31_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_15 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_16  (
    .i0(inst_doa_i32_001),
    .i1(inst_doa_i33_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_16 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_17  (
    .i0(inst_doa_i34_001),
    .i1(inst_doa_i35_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_17 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_18  (
    .i0(inst_doa_i36_001),
    .i1(inst_doa_i37_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_18 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_19  (
    .i0(inst_doa_i38_001),
    .i1(inst_doa_i39_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_19 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_2  (
    .i0(inst_doa_i4_001),
    .i1(inst_doa_i5_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_2 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_20  (
    .i0(inst_doa_i40_001),
    .i1(inst_doa_i41_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_20 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_21  (
    .i0(inst_doa_i42_001),
    .i1(inst_doa_i43_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_21 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_22  (
    .i0(inst_doa_i44_001),
    .i1(inst_doa_i45_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_22 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_23  (
    .i0(inst_doa_i46_001),
    .i1(inst_doa_i47_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_23 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_24  (
    .i0(inst_doa_i48_001),
    .i1(inst_doa_i49_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_24 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_25  (
    .i0(inst_doa_i50_001),
    .i1(inst_doa_i51_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_25 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_26  (
    .i0(inst_doa_i52_001),
    .i1(inst_doa_i53_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_26 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_27  (
    .i0(inst_doa_i54_001),
    .i1(inst_doa_i55_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_27 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_28  (
    .i0(inst_doa_i56_001),
    .i1(inst_doa_i57_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_28 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_29  (
    .i0(inst_doa_i58_001),
    .i1(inst_doa_i59_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_29 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_3  (
    .i0(inst_doa_i6_001),
    .i1(inst_doa_i7_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_3 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_30  (
    .i0(inst_doa_i60_001),
    .i1(inst_doa_i61_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_30 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_31  (
    .i0(inst_doa_i62_001),
    .i1(inst_doa_i63_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_31 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_4  (
    .i0(inst_doa_i8_001),
    .i1(inst_doa_i9_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_4 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_5  (
    .i0(inst_doa_i10_001),
    .i1(inst_doa_i11_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_5 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_6  (
    .i0(inst_doa_i12_001),
    .i1(inst_doa_i13_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_6 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_7  (
    .i0(inst_doa_i14_001),
    .i1(inst_doa_i15_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_7 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_8  (
    .i0(inst_doa_i16_001),
    .i1(inst_doa_i17_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_8 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_9  (
    .i0(inst_doa_i18_001),
    .i1(inst_doa_i19_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_9 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b1/B0_0 ),
    .i1(\inst_doa_mux_b1/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_0 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b1/B0_2 ),
    .i1(\inst_doa_mux_b1/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_1 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_10  (
    .i0(\inst_doa_mux_b1/B0_20 ),
    .i1(\inst_doa_mux_b1/B0_21 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_10 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_11  (
    .i0(\inst_doa_mux_b1/B0_22 ),
    .i1(\inst_doa_mux_b1/B0_23 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_11 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_12  (
    .i0(\inst_doa_mux_b1/B0_24 ),
    .i1(\inst_doa_mux_b1/B0_25 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_12 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_13  (
    .i0(\inst_doa_mux_b1/B0_26 ),
    .i1(\inst_doa_mux_b1/B0_27 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_13 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_14  (
    .i0(\inst_doa_mux_b1/B0_28 ),
    .i1(\inst_doa_mux_b1/B0_29 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_14 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_15  (
    .i0(\inst_doa_mux_b1/B0_30 ),
    .i1(\inst_doa_mux_b1/B0_31 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_15 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_2  (
    .i0(\inst_doa_mux_b1/B0_4 ),
    .i1(\inst_doa_mux_b1/B0_5 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_2 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_3  (
    .i0(\inst_doa_mux_b1/B0_6 ),
    .i1(\inst_doa_mux_b1/B0_7 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_3 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_4  (
    .i0(\inst_doa_mux_b1/B0_8 ),
    .i1(\inst_doa_mux_b1/B0_9 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_4 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_5  (
    .i0(\inst_doa_mux_b1/B0_10 ),
    .i1(\inst_doa_mux_b1/B0_11 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_5 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_6  (
    .i0(\inst_doa_mux_b1/B0_12 ),
    .i1(\inst_doa_mux_b1/B0_13 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_6 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_7  (
    .i0(\inst_doa_mux_b1/B0_14 ),
    .i1(\inst_doa_mux_b1/B0_15 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_7 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_8  (
    .i0(\inst_doa_mux_b1/B0_16 ),
    .i1(\inst_doa_mux_b1/B0_17 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_8 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_9  (
    .i0(\inst_doa_mux_b1/B0_18 ),
    .i1(\inst_doa_mux_b1/B0_19 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_9 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b1/B1_0 ),
    .i1(\inst_doa_mux_b1/B1_1 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b1/B2_0 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_2_1  (
    .i0(\inst_doa_mux_b1/B1_2 ),
    .i1(\inst_doa_mux_b1/B1_3 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b1/B2_1 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_2_2  (
    .i0(\inst_doa_mux_b1/B1_4 ),
    .i1(\inst_doa_mux_b1/B1_5 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b1/B2_2 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_2_3  (
    .i0(\inst_doa_mux_b1/B1_6 ),
    .i1(\inst_doa_mux_b1/B1_7 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b1/B2_3 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_2_4  (
    .i0(\inst_doa_mux_b1/B1_8 ),
    .i1(\inst_doa_mux_b1/B1_9 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b1/B2_4 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_2_5  (
    .i0(\inst_doa_mux_b1/B1_10 ),
    .i1(\inst_doa_mux_b1/B1_11 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b1/B2_5 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_2_6  (
    .i0(\inst_doa_mux_b1/B1_12 ),
    .i1(\inst_doa_mux_b1/B1_13 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b1/B2_6 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_2_7  (
    .i0(\inst_doa_mux_b1/B1_14 ),
    .i1(\inst_doa_mux_b1/B1_15 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b1/B2_7 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_3_0  (
    .i0(\inst_doa_mux_b1/B2_0 ),
    .i1(\inst_doa_mux_b1/B2_1 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b1/B3_0 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_3_1  (
    .i0(\inst_doa_mux_b1/B2_2 ),
    .i1(\inst_doa_mux_b1/B2_3 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b1/B3_1 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_3_2  (
    .i0(\inst_doa_mux_b1/B2_4 ),
    .i1(\inst_doa_mux_b1/B2_5 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b1/B3_2 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_3_3  (
    .i0(\inst_doa_mux_b1/B2_6 ),
    .i1(\inst_doa_mux_b1/B2_7 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b1/B3_3 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_4_0  (
    .i0(\inst_doa_mux_b1/B3_0 ),
    .i1(\inst_doa_mux_b1/B3_1 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b1/B4_0 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_4_1  (
    .i0(\inst_doa_mux_b1/B3_2 ),
    .i1(\inst_doa_mux_b1/B3_3 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b1/B4_1 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_5_0  (
    .i0(\inst_doa_mux_b1/B4_0 ),
    .i1(\inst_doa_mux_b1/B4_1 ),
    .sel(addra_piped[5]),
    .o(doa[1]));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_3_0  (
    .i0(inst_doa_i0_010),
    .i1(inst_doa_i8_010),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b10/B3_0 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_3_1  (
    .i0(inst_doa_i16_010),
    .i1(inst_doa_i24_010),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b10/B3_1 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_3_2  (
    .i0(inst_doa_i32_010),
    .i1(inst_doa_i40_010),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b10/B3_2 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_3_3  (
    .i0(inst_doa_i48_010),
    .i1(inst_doa_i56_010),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b10/B3_3 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_4_0  (
    .i0(\inst_doa_mux_b10/B3_0 ),
    .i1(\inst_doa_mux_b10/B3_1 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b10/B4_0 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_4_1  (
    .i0(\inst_doa_mux_b10/B3_2 ),
    .i1(\inst_doa_mux_b10/B3_3 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b10/B4_1 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_5_0  (
    .i0(\inst_doa_mux_b10/B4_0 ),
    .i1(\inst_doa_mux_b10/B4_1 ),
    .sel(addra_piped[5]),
    .o(doa[10]));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_3_0  (
    .i0(inst_doa_i0_010),
    .i1(inst_doa_i8_011),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b11/B3_0 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_3_1  (
    .i0(inst_doa_i16_011),
    .i1(inst_doa_i24_010),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b11/B3_1 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_3_2  (
    .i0(inst_doa_i32_010),
    .i1(inst_doa_i40_011),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b11/B3_2 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_3_3  (
    .i0(inst_doa_i48_011),
    .i1(inst_doa_i56_010),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b11/B3_3 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_4_0  (
    .i0(\inst_doa_mux_b11/B3_0 ),
    .i1(\inst_doa_mux_b11/B3_1 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b11/B4_0 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_4_1  (
    .i0(\inst_doa_mux_b11/B3_2 ),
    .i1(\inst_doa_mux_b11/B3_3 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b11/B4_1 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_5_0  (
    .i0(\inst_doa_mux_b11/B4_0 ),
    .i1(\inst_doa_mux_b11/B4_1 ),
    .sel(addra_piped[5]),
    .o(doa[11]));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_0  (
    .i0(inst_doa_i0_002),
    .i1(inst_doa_i1_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_0 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_1  (
    .i0(inst_doa_i2_002),
    .i1(inst_doa_i3_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_1 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_10  (
    .i0(inst_doa_i20_002),
    .i1(inst_doa_i21_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_10 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_11  (
    .i0(inst_doa_i22_002),
    .i1(inst_doa_i23_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_11 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_12  (
    .i0(inst_doa_i24_002),
    .i1(inst_doa_i25_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_12 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_13  (
    .i0(inst_doa_i26_002),
    .i1(inst_doa_i27_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_13 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_14  (
    .i0(inst_doa_i28_002),
    .i1(inst_doa_i29_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_14 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_15  (
    .i0(inst_doa_i30_002),
    .i1(inst_doa_i31_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_15 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_16  (
    .i0(inst_doa_i32_002),
    .i1(inst_doa_i33_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_16 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_17  (
    .i0(inst_doa_i34_002),
    .i1(inst_doa_i35_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_17 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_18  (
    .i0(inst_doa_i36_002),
    .i1(inst_doa_i37_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_18 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_19  (
    .i0(inst_doa_i38_002),
    .i1(inst_doa_i39_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_19 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_2  (
    .i0(inst_doa_i4_002),
    .i1(inst_doa_i5_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_2 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_20  (
    .i0(inst_doa_i40_002),
    .i1(inst_doa_i41_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_20 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_21  (
    .i0(inst_doa_i42_002),
    .i1(inst_doa_i43_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_21 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_22  (
    .i0(inst_doa_i44_002),
    .i1(inst_doa_i45_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_22 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_23  (
    .i0(inst_doa_i46_002),
    .i1(inst_doa_i47_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_23 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_24  (
    .i0(inst_doa_i48_002),
    .i1(inst_doa_i49_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_24 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_25  (
    .i0(inst_doa_i50_002),
    .i1(inst_doa_i51_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_25 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_26  (
    .i0(inst_doa_i52_002),
    .i1(inst_doa_i53_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_26 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_27  (
    .i0(inst_doa_i54_002),
    .i1(inst_doa_i55_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_27 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_28  (
    .i0(inst_doa_i56_002),
    .i1(inst_doa_i57_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_28 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_29  (
    .i0(inst_doa_i58_002),
    .i1(inst_doa_i59_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_29 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_3  (
    .i0(inst_doa_i6_002),
    .i1(inst_doa_i7_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_3 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_30  (
    .i0(inst_doa_i60_002),
    .i1(inst_doa_i61_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_30 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_31  (
    .i0(inst_doa_i62_002),
    .i1(inst_doa_i63_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_31 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_4  (
    .i0(inst_doa_i8_002),
    .i1(inst_doa_i9_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_4 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_5  (
    .i0(inst_doa_i10_002),
    .i1(inst_doa_i11_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_5 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_6  (
    .i0(inst_doa_i12_002),
    .i1(inst_doa_i13_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_6 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_7  (
    .i0(inst_doa_i14_002),
    .i1(inst_doa_i15_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_7 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_8  (
    .i0(inst_doa_i16_002),
    .i1(inst_doa_i17_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_8 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_9  (
    .i0(inst_doa_i18_002),
    .i1(inst_doa_i19_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_9 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b2/B0_0 ),
    .i1(\inst_doa_mux_b2/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_0 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b2/B0_2 ),
    .i1(\inst_doa_mux_b2/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_1 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_10  (
    .i0(\inst_doa_mux_b2/B0_20 ),
    .i1(\inst_doa_mux_b2/B0_21 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_10 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_11  (
    .i0(\inst_doa_mux_b2/B0_22 ),
    .i1(\inst_doa_mux_b2/B0_23 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_11 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_12  (
    .i0(\inst_doa_mux_b2/B0_24 ),
    .i1(\inst_doa_mux_b2/B0_25 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_12 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_13  (
    .i0(\inst_doa_mux_b2/B0_26 ),
    .i1(\inst_doa_mux_b2/B0_27 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_13 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_14  (
    .i0(\inst_doa_mux_b2/B0_28 ),
    .i1(\inst_doa_mux_b2/B0_29 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_14 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_15  (
    .i0(\inst_doa_mux_b2/B0_30 ),
    .i1(\inst_doa_mux_b2/B0_31 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_15 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_2  (
    .i0(\inst_doa_mux_b2/B0_4 ),
    .i1(\inst_doa_mux_b2/B0_5 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_2 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_3  (
    .i0(\inst_doa_mux_b2/B0_6 ),
    .i1(\inst_doa_mux_b2/B0_7 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_3 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_4  (
    .i0(\inst_doa_mux_b2/B0_8 ),
    .i1(\inst_doa_mux_b2/B0_9 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_4 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_5  (
    .i0(\inst_doa_mux_b2/B0_10 ),
    .i1(\inst_doa_mux_b2/B0_11 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_5 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_6  (
    .i0(\inst_doa_mux_b2/B0_12 ),
    .i1(\inst_doa_mux_b2/B0_13 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_6 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_7  (
    .i0(\inst_doa_mux_b2/B0_14 ),
    .i1(\inst_doa_mux_b2/B0_15 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_7 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_8  (
    .i0(\inst_doa_mux_b2/B0_16 ),
    .i1(\inst_doa_mux_b2/B0_17 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_8 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_9  (
    .i0(\inst_doa_mux_b2/B0_18 ),
    .i1(\inst_doa_mux_b2/B0_19 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_9 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b2/B1_0 ),
    .i1(\inst_doa_mux_b2/B1_1 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b2/B2_0 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_2_1  (
    .i0(\inst_doa_mux_b2/B1_2 ),
    .i1(\inst_doa_mux_b2/B1_3 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b2/B2_1 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_2_2  (
    .i0(\inst_doa_mux_b2/B1_4 ),
    .i1(\inst_doa_mux_b2/B1_5 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b2/B2_2 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_2_3  (
    .i0(\inst_doa_mux_b2/B1_6 ),
    .i1(\inst_doa_mux_b2/B1_7 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b2/B2_3 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_2_4  (
    .i0(\inst_doa_mux_b2/B1_8 ),
    .i1(\inst_doa_mux_b2/B1_9 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b2/B2_4 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_2_5  (
    .i0(\inst_doa_mux_b2/B1_10 ),
    .i1(\inst_doa_mux_b2/B1_11 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b2/B2_5 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_2_6  (
    .i0(\inst_doa_mux_b2/B1_12 ),
    .i1(\inst_doa_mux_b2/B1_13 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b2/B2_6 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_2_7  (
    .i0(\inst_doa_mux_b2/B1_14 ),
    .i1(\inst_doa_mux_b2/B1_15 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b2/B2_7 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_3_0  (
    .i0(\inst_doa_mux_b2/B2_0 ),
    .i1(\inst_doa_mux_b2/B2_1 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b2/B3_0 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_3_1  (
    .i0(\inst_doa_mux_b2/B2_2 ),
    .i1(\inst_doa_mux_b2/B2_3 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b2/B3_1 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_3_2  (
    .i0(\inst_doa_mux_b2/B2_4 ),
    .i1(\inst_doa_mux_b2/B2_5 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b2/B3_2 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_3_3  (
    .i0(\inst_doa_mux_b2/B2_6 ),
    .i1(\inst_doa_mux_b2/B2_7 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b2/B3_3 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_4_0  (
    .i0(\inst_doa_mux_b2/B3_0 ),
    .i1(\inst_doa_mux_b2/B3_1 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b2/B4_0 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_4_1  (
    .i0(\inst_doa_mux_b2/B3_2 ),
    .i1(\inst_doa_mux_b2/B3_3 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b2/B4_1 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_5_0  (
    .i0(\inst_doa_mux_b2/B4_0 ),
    .i1(\inst_doa_mux_b2/B4_1 ),
    .sel(addra_piped[5]),
    .o(doa[2]));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_0  (
    .i0(inst_doa_i0_003),
    .i1(inst_doa_i1_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_0 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_1  (
    .i0(inst_doa_i2_003),
    .i1(inst_doa_i3_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_1 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_10  (
    .i0(inst_doa_i20_003),
    .i1(inst_doa_i21_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_10 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_11  (
    .i0(inst_doa_i22_003),
    .i1(inst_doa_i23_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_11 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_12  (
    .i0(inst_doa_i24_003),
    .i1(inst_doa_i25_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_12 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_13  (
    .i0(inst_doa_i26_003),
    .i1(inst_doa_i27_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_13 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_14  (
    .i0(inst_doa_i28_003),
    .i1(inst_doa_i29_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_14 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_15  (
    .i0(inst_doa_i30_003),
    .i1(inst_doa_i31_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_15 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_16  (
    .i0(inst_doa_i32_003),
    .i1(inst_doa_i33_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_16 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_17  (
    .i0(inst_doa_i34_003),
    .i1(inst_doa_i35_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_17 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_18  (
    .i0(inst_doa_i36_003),
    .i1(inst_doa_i37_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_18 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_19  (
    .i0(inst_doa_i38_003),
    .i1(inst_doa_i39_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_19 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_2  (
    .i0(inst_doa_i4_003),
    .i1(inst_doa_i5_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_2 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_20  (
    .i0(inst_doa_i40_003),
    .i1(inst_doa_i41_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_20 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_21  (
    .i0(inst_doa_i42_003),
    .i1(inst_doa_i43_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_21 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_22  (
    .i0(inst_doa_i44_003),
    .i1(inst_doa_i45_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_22 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_23  (
    .i0(inst_doa_i46_003),
    .i1(inst_doa_i47_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_23 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_24  (
    .i0(inst_doa_i48_003),
    .i1(inst_doa_i49_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_24 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_25  (
    .i0(inst_doa_i50_003),
    .i1(inst_doa_i51_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_25 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_26  (
    .i0(inst_doa_i52_003),
    .i1(inst_doa_i53_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_26 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_27  (
    .i0(inst_doa_i54_003),
    .i1(inst_doa_i55_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_27 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_28  (
    .i0(inst_doa_i56_003),
    .i1(inst_doa_i57_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_28 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_29  (
    .i0(inst_doa_i58_003),
    .i1(inst_doa_i59_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_29 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_3  (
    .i0(inst_doa_i6_003),
    .i1(inst_doa_i7_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_3 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_30  (
    .i0(inst_doa_i60_003),
    .i1(inst_doa_i61_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_30 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_31  (
    .i0(inst_doa_i62_003),
    .i1(inst_doa_i63_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_31 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_4  (
    .i0(inst_doa_i8_003),
    .i1(inst_doa_i9_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_4 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_5  (
    .i0(inst_doa_i10_003),
    .i1(inst_doa_i11_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_5 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_6  (
    .i0(inst_doa_i12_003),
    .i1(inst_doa_i13_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_6 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_7  (
    .i0(inst_doa_i14_003),
    .i1(inst_doa_i15_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_7 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_8  (
    .i0(inst_doa_i16_003),
    .i1(inst_doa_i17_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_8 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_9  (
    .i0(inst_doa_i18_003),
    .i1(inst_doa_i19_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_9 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b3/B0_0 ),
    .i1(\inst_doa_mux_b3/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_0 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b3/B0_2 ),
    .i1(\inst_doa_mux_b3/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_1 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_10  (
    .i0(\inst_doa_mux_b3/B0_20 ),
    .i1(\inst_doa_mux_b3/B0_21 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_10 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_11  (
    .i0(\inst_doa_mux_b3/B0_22 ),
    .i1(\inst_doa_mux_b3/B0_23 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_11 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_12  (
    .i0(\inst_doa_mux_b3/B0_24 ),
    .i1(\inst_doa_mux_b3/B0_25 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_12 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_13  (
    .i0(\inst_doa_mux_b3/B0_26 ),
    .i1(\inst_doa_mux_b3/B0_27 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_13 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_14  (
    .i0(\inst_doa_mux_b3/B0_28 ),
    .i1(\inst_doa_mux_b3/B0_29 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_14 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_15  (
    .i0(\inst_doa_mux_b3/B0_30 ),
    .i1(\inst_doa_mux_b3/B0_31 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_15 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_2  (
    .i0(\inst_doa_mux_b3/B0_4 ),
    .i1(\inst_doa_mux_b3/B0_5 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_2 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_3  (
    .i0(\inst_doa_mux_b3/B0_6 ),
    .i1(\inst_doa_mux_b3/B0_7 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_3 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_4  (
    .i0(\inst_doa_mux_b3/B0_8 ),
    .i1(\inst_doa_mux_b3/B0_9 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_4 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_5  (
    .i0(\inst_doa_mux_b3/B0_10 ),
    .i1(\inst_doa_mux_b3/B0_11 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_5 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_6  (
    .i0(\inst_doa_mux_b3/B0_12 ),
    .i1(\inst_doa_mux_b3/B0_13 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_6 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_7  (
    .i0(\inst_doa_mux_b3/B0_14 ),
    .i1(\inst_doa_mux_b3/B0_15 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_7 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_8  (
    .i0(\inst_doa_mux_b3/B0_16 ),
    .i1(\inst_doa_mux_b3/B0_17 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_8 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_9  (
    .i0(\inst_doa_mux_b3/B0_18 ),
    .i1(\inst_doa_mux_b3/B0_19 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_9 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b3/B1_0 ),
    .i1(\inst_doa_mux_b3/B1_1 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b3/B2_0 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_2_1  (
    .i0(\inst_doa_mux_b3/B1_2 ),
    .i1(\inst_doa_mux_b3/B1_3 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b3/B2_1 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_2_2  (
    .i0(\inst_doa_mux_b3/B1_4 ),
    .i1(\inst_doa_mux_b3/B1_5 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b3/B2_2 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_2_3  (
    .i0(\inst_doa_mux_b3/B1_6 ),
    .i1(\inst_doa_mux_b3/B1_7 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b3/B2_3 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_2_4  (
    .i0(\inst_doa_mux_b3/B1_8 ),
    .i1(\inst_doa_mux_b3/B1_9 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b3/B2_4 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_2_5  (
    .i0(\inst_doa_mux_b3/B1_10 ),
    .i1(\inst_doa_mux_b3/B1_11 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b3/B2_5 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_2_6  (
    .i0(\inst_doa_mux_b3/B1_12 ),
    .i1(\inst_doa_mux_b3/B1_13 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b3/B2_6 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_2_7  (
    .i0(\inst_doa_mux_b3/B1_14 ),
    .i1(\inst_doa_mux_b3/B1_15 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b3/B2_7 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_3_0  (
    .i0(\inst_doa_mux_b3/B2_0 ),
    .i1(\inst_doa_mux_b3/B2_1 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b3/B3_0 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_3_1  (
    .i0(\inst_doa_mux_b3/B2_2 ),
    .i1(\inst_doa_mux_b3/B2_3 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b3/B3_1 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_3_2  (
    .i0(\inst_doa_mux_b3/B2_4 ),
    .i1(\inst_doa_mux_b3/B2_5 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b3/B3_2 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_3_3  (
    .i0(\inst_doa_mux_b3/B2_6 ),
    .i1(\inst_doa_mux_b3/B2_7 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b3/B3_3 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_4_0  (
    .i0(\inst_doa_mux_b3/B3_0 ),
    .i1(\inst_doa_mux_b3/B3_1 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b3/B4_0 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_4_1  (
    .i0(\inst_doa_mux_b3/B3_2 ),
    .i1(\inst_doa_mux_b3/B3_3 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b3/B4_1 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_5_0  (
    .i0(\inst_doa_mux_b3/B4_0 ),
    .i1(\inst_doa_mux_b3/B4_1 ),
    .sel(addra_piped[5]),
    .o(doa[3]));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_0  (
    .i0(inst_doa_i0_004),
    .i1(inst_doa_i1_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_0 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_1  (
    .i0(inst_doa_i2_004),
    .i1(inst_doa_i3_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_1 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_10  (
    .i0(inst_doa_i20_004),
    .i1(inst_doa_i21_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_10 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_11  (
    .i0(inst_doa_i22_004),
    .i1(inst_doa_i23_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_11 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_12  (
    .i0(inst_doa_i24_004),
    .i1(inst_doa_i25_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_12 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_13  (
    .i0(inst_doa_i26_004),
    .i1(inst_doa_i27_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_13 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_14  (
    .i0(inst_doa_i28_004),
    .i1(inst_doa_i29_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_14 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_15  (
    .i0(inst_doa_i30_004),
    .i1(inst_doa_i31_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_15 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_16  (
    .i0(inst_doa_i32_004),
    .i1(inst_doa_i33_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_16 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_17  (
    .i0(inst_doa_i34_004),
    .i1(inst_doa_i35_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_17 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_18  (
    .i0(inst_doa_i36_004),
    .i1(inst_doa_i37_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_18 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_19  (
    .i0(inst_doa_i38_004),
    .i1(inst_doa_i39_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_19 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_2  (
    .i0(inst_doa_i4_004),
    .i1(inst_doa_i5_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_2 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_20  (
    .i0(inst_doa_i40_004),
    .i1(inst_doa_i41_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_20 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_21  (
    .i0(inst_doa_i42_004),
    .i1(inst_doa_i43_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_21 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_22  (
    .i0(inst_doa_i44_004),
    .i1(inst_doa_i45_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_22 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_23  (
    .i0(inst_doa_i46_004),
    .i1(inst_doa_i47_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_23 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_24  (
    .i0(inst_doa_i48_004),
    .i1(inst_doa_i49_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_24 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_25  (
    .i0(inst_doa_i50_004),
    .i1(inst_doa_i51_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_25 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_26  (
    .i0(inst_doa_i52_004),
    .i1(inst_doa_i53_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_26 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_27  (
    .i0(inst_doa_i54_004),
    .i1(inst_doa_i55_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_27 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_28  (
    .i0(inst_doa_i56_004),
    .i1(inst_doa_i57_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_28 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_29  (
    .i0(inst_doa_i58_004),
    .i1(inst_doa_i59_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_29 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_3  (
    .i0(inst_doa_i6_004),
    .i1(inst_doa_i7_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_3 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_30  (
    .i0(inst_doa_i60_004),
    .i1(inst_doa_i61_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_30 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_31  (
    .i0(inst_doa_i62_004),
    .i1(inst_doa_i63_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_31 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_4  (
    .i0(inst_doa_i8_004),
    .i1(inst_doa_i9_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_4 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_5  (
    .i0(inst_doa_i10_004),
    .i1(inst_doa_i11_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_5 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_6  (
    .i0(inst_doa_i12_004),
    .i1(inst_doa_i13_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_6 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_7  (
    .i0(inst_doa_i14_004),
    .i1(inst_doa_i15_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_7 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_8  (
    .i0(inst_doa_i16_004),
    .i1(inst_doa_i17_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_8 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_9  (
    .i0(inst_doa_i18_004),
    .i1(inst_doa_i19_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_9 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b4/B0_0 ),
    .i1(\inst_doa_mux_b4/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_0 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b4/B0_2 ),
    .i1(\inst_doa_mux_b4/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_1 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_10  (
    .i0(\inst_doa_mux_b4/B0_20 ),
    .i1(\inst_doa_mux_b4/B0_21 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_10 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_11  (
    .i0(\inst_doa_mux_b4/B0_22 ),
    .i1(\inst_doa_mux_b4/B0_23 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_11 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_12  (
    .i0(\inst_doa_mux_b4/B0_24 ),
    .i1(\inst_doa_mux_b4/B0_25 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_12 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_13  (
    .i0(\inst_doa_mux_b4/B0_26 ),
    .i1(\inst_doa_mux_b4/B0_27 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_13 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_14  (
    .i0(\inst_doa_mux_b4/B0_28 ),
    .i1(\inst_doa_mux_b4/B0_29 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_14 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_15  (
    .i0(\inst_doa_mux_b4/B0_30 ),
    .i1(\inst_doa_mux_b4/B0_31 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_15 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_2  (
    .i0(\inst_doa_mux_b4/B0_4 ),
    .i1(\inst_doa_mux_b4/B0_5 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_2 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_3  (
    .i0(\inst_doa_mux_b4/B0_6 ),
    .i1(\inst_doa_mux_b4/B0_7 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_3 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_4  (
    .i0(\inst_doa_mux_b4/B0_8 ),
    .i1(\inst_doa_mux_b4/B0_9 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_4 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_5  (
    .i0(\inst_doa_mux_b4/B0_10 ),
    .i1(\inst_doa_mux_b4/B0_11 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_5 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_6  (
    .i0(\inst_doa_mux_b4/B0_12 ),
    .i1(\inst_doa_mux_b4/B0_13 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_6 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_7  (
    .i0(\inst_doa_mux_b4/B0_14 ),
    .i1(\inst_doa_mux_b4/B0_15 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_7 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_8  (
    .i0(\inst_doa_mux_b4/B0_16 ),
    .i1(\inst_doa_mux_b4/B0_17 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_8 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_9  (
    .i0(\inst_doa_mux_b4/B0_18 ),
    .i1(\inst_doa_mux_b4/B0_19 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_9 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b4/B1_0 ),
    .i1(\inst_doa_mux_b4/B1_1 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b4/B2_0 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_2_1  (
    .i0(\inst_doa_mux_b4/B1_2 ),
    .i1(\inst_doa_mux_b4/B1_3 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b4/B2_1 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_2_2  (
    .i0(\inst_doa_mux_b4/B1_4 ),
    .i1(\inst_doa_mux_b4/B1_5 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b4/B2_2 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_2_3  (
    .i0(\inst_doa_mux_b4/B1_6 ),
    .i1(\inst_doa_mux_b4/B1_7 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b4/B2_3 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_2_4  (
    .i0(\inst_doa_mux_b4/B1_8 ),
    .i1(\inst_doa_mux_b4/B1_9 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b4/B2_4 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_2_5  (
    .i0(\inst_doa_mux_b4/B1_10 ),
    .i1(\inst_doa_mux_b4/B1_11 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b4/B2_5 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_2_6  (
    .i0(\inst_doa_mux_b4/B1_12 ),
    .i1(\inst_doa_mux_b4/B1_13 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b4/B2_6 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_2_7  (
    .i0(\inst_doa_mux_b4/B1_14 ),
    .i1(\inst_doa_mux_b4/B1_15 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b4/B2_7 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_3_0  (
    .i0(\inst_doa_mux_b4/B2_0 ),
    .i1(\inst_doa_mux_b4/B2_1 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b4/B3_0 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_3_1  (
    .i0(\inst_doa_mux_b4/B2_2 ),
    .i1(\inst_doa_mux_b4/B2_3 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b4/B3_1 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_3_2  (
    .i0(\inst_doa_mux_b4/B2_4 ),
    .i1(\inst_doa_mux_b4/B2_5 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b4/B3_2 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_3_3  (
    .i0(\inst_doa_mux_b4/B2_6 ),
    .i1(\inst_doa_mux_b4/B2_7 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b4/B3_3 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_4_0  (
    .i0(\inst_doa_mux_b4/B3_0 ),
    .i1(\inst_doa_mux_b4/B3_1 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b4/B4_0 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_4_1  (
    .i0(\inst_doa_mux_b4/B3_2 ),
    .i1(\inst_doa_mux_b4/B3_3 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b4/B4_1 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_5_0  (
    .i0(\inst_doa_mux_b4/B4_0 ),
    .i1(\inst_doa_mux_b4/B4_1 ),
    .sel(addra_piped[5]),
    .o(doa[4]));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_0  (
    .i0(inst_doa_i0_005),
    .i1(inst_doa_i1_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_0 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_1  (
    .i0(inst_doa_i2_005),
    .i1(inst_doa_i3_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_1 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_10  (
    .i0(inst_doa_i20_005),
    .i1(inst_doa_i21_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_10 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_11  (
    .i0(inst_doa_i22_005),
    .i1(inst_doa_i23_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_11 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_12  (
    .i0(inst_doa_i24_005),
    .i1(inst_doa_i25_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_12 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_13  (
    .i0(inst_doa_i26_005),
    .i1(inst_doa_i27_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_13 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_14  (
    .i0(inst_doa_i28_005),
    .i1(inst_doa_i29_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_14 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_15  (
    .i0(inst_doa_i30_005),
    .i1(inst_doa_i31_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_15 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_16  (
    .i0(inst_doa_i32_005),
    .i1(inst_doa_i33_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_16 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_17  (
    .i0(inst_doa_i34_005),
    .i1(inst_doa_i35_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_17 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_18  (
    .i0(inst_doa_i36_005),
    .i1(inst_doa_i37_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_18 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_19  (
    .i0(inst_doa_i38_005),
    .i1(inst_doa_i39_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_19 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_2  (
    .i0(inst_doa_i4_005),
    .i1(inst_doa_i5_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_2 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_20  (
    .i0(inst_doa_i40_005),
    .i1(inst_doa_i41_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_20 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_21  (
    .i0(inst_doa_i42_005),
    .i1(inst_doa_i43_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_21 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_22  (
    .i0(inst_doa_i44_005),
    .i1(inst_doa_i45_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_22 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_23  (
    .i0(inst_doa_i46_005),
    .i1(inst_doa_i47_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_23 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_24  (
    .i0(inst_doa_i48_005),
    .i1(inst_doa_i49_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_24 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_25  (
    .i0(inst_doa_i50_005),
    .i1(inst_doa_i51_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_25 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_26  (
    .i0(inst_doa_i52_005),
    .i1(inst_doa_i53_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_26 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_27  (
    .i0(inst_doa_i54_005),
    .i1(inst_doa_i55_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_27 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_28  (
    .i0(inst_doa_i56_005),
    .i1(inst_doa_i57_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_28 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_29  (
    .i0(inst_doa_i58_005),
    .i1(inst_doa_i59_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_29 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_3  (
    .i0(inst_doa_i6_005),
    .i1(inst_doa_i7_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_3 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_30  (
    .i0(inst_doa_i60_005),
    .i1(inst_doa_i61_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_30 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_31  (
    .i0(inst_doa_i62_005),
    .i1(inst_doa_i63_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_31 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_4  (
    .i0(inst_doa_i8_005),
    .i1(inst_doa_i9_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_4 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_5  (
    .i0(inst_doa_i10_005),
    .i1(inst_doa_i11_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_5 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_6  (
    .i0(inst_doa_i12_005),
    .i1(inst_doa_i13_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_6 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_7  (
    .i0(inst_doa_i14_005),
    .i1(inst_doa_i15_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_7 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_8  (
    .i0(inst_doa_i16_005),
    .i1(inst_doa_i17_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_8 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_9  (
    .i0(inst_doa_i18_005),
    .i1(inst_doa_i19_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_9 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b5/B0_0 ),
    .i1(\inst_doa_mux_b5/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_0 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b5/B0_2 ),
    .i1(\inst_doa_mux_b5/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_1 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_10  (
    .i0(\inst_doa_mux_b5/B0_20 ),
    .i1(\inst_doa_mux_b5/B0_21 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_10 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_11  (
    .i0(\inst_doa_mux_b5/B0_22 ),
    .i1(\inst_doa_mux_b5/B0_23 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_11 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_12  (
    .i0(\inst_doa_mux_b5/B0_24 ),
    .i1(\inst_doa_mux_b5/B0_25 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_12 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_13  (
    .i0(\inst_doa_mux_b5/B0_26 ),
    .i1(\inst_doa_mux_b5/B0_27 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_13 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_14  (
    .i0(\inst_doa_mux_b5/B0_28 ),
    .i1(\inst_doa_mux_b5/B0_29 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_14 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_15  (
    .i0(\inst_doa_mux_b5/B0_30 ),
    .i1(\inst_doa_mux_b5/B0_31 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_15 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_2  (
    .i0(\inst_doa_mux_b5/B0_4 ),
    .i1(\inst_doa_mux_b5/B0_5 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_2 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_3  (
    .i0(\inst_doa_mux_b5/B0_6 ),
    .i1(\inst_doa_mux_b5/B0_7 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_3 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_4  (
    .i0(\inst_doa_mux_b5/B0_8 ),
    .i1(\inst_doa_mux_b5/B0_9 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_4 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_5  (
    .i0(\inst_doa_mux_b5/B0_10 ),
    .i1(\inst_doa_mux_b5/B0_11 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_5 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_6  (
    .i0(\inst_doa_mux_b5/B0_12 ),
    .i1(\inst_doa_mux_b5/B0_13 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_6 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_7  (
    .i0(\inst_doa_mux_b5/B0_14 ),
    .i1(\inst_doa_mux_b5/B0_15 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_7 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_8  (
    .i0(\inst_doa_mux_b5/B0_16 ),
    .i1(\inst_doa_mux_b5/B0_17 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_8 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_9  (
    .i0(\inst_doa_mux_b5/B0_18 ),
    .i1(\inst_doa_mux_b5/B0_19 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_9 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b5/B1_0 ),
    .i1(\inst_doa_mux_b5/B1_1 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b5/B2_0 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_2_1  (
    .i0(\inst_doa_mux_b5/B1_2 ),
    .i1(\inst_doa_mux_b5/B1_3 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b5/B2_1 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_2_2  (
    .i0(\inst_doa_mux_b5/B1_4 ),
    .i1(\inst_doa_mux_b5/B1_5 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b5/B2_2 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_2_3  (
    .i0(\inst_doa_mux_b5/B1_6 ),
    .i1(\inst_doa_mux_b5/B1_7 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b5/B2_3 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_2_4  (
    .i0(\inst_doa_mux_b5/B1_8 ),
    .i1(\inst_doa_mux_b5/B1_9 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b5/B2_4 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_2_5  (
    .i0(\inst_doa_mux_b5/B1_10 ),
    .i1(\inst_doa_mux_b5/B1_11 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b5/B2_5 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_2_6  (
    .i0(\inst_doa_mux_b5/B1_12 ),
    .i1(\inst_doa_mux_b5/B1_13 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b5/B2_6 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_2_7  (
    .i0(\inst_doa_mux_b5/B1_14 ),
    .i1(\inst_doa_mux_b5/B1_15 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b5/B2_7 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_3_0  (
    .i0(\inst_doa_mux_b5/B2_0 ),
    .i1(\inst_doa_mux_b5/B2_1 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b5/B3_0 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_3_1  (
    .i0(\inst_doa_mux_b5/B2_2 ),
    .i1(\inst_doa_mux_b5/B2_3 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b5/B3_1 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_3_2  (
    .i0(\inst_doa_mux_b5/B2_4 ),
    .i1(\inst_doa_mux_b5/B2_5 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b5/B3_2 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_3_3  (
    .i0(\inst_doa_mux_b5/B2_6 ),
    .i1(\inst_doa_mux_b5/B2_7 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b5/B3_3 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_4_0  (
    .i0(\inst_doa_mux_b5/B3_0 ),
    .i1(\inst_doa_mux_b5/B3_1 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b5/B4_0 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_4_1  (
    .i0(\inst_doa_mux_b5/B3_2 ),
    .i1(\inst_doa_mux_b5/B3_3 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b5/B4_1 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_5_0  (
    .i0(\inst_doa_mux_b5/B4_0 ),
    .i1(\inst_doa_mux_b5/B4_1 ),
    .sel(addra_piped[5]),
    .o(doa[5]));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_0  (
    .i0(inst_doa_i0_006),
    .i1(inst_doa_i1_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_0 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_1  (
    .i0(inst_doa_i2_006),
    .i1(inst_doa_i3_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_1 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_10  (
    .i0(inst_doa_i20_006),
    .i1(inst_doa_i21_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_10 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_11  (
    .i0(inst_doa_i22_006),
    .i1(inst_doa_i23_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_11 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_12  (
    .i0(inst_doa_i24_006),
    .i1(inst_doa_i25_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_12 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_13  (
    .i0(inst_doa_i26_006),
    .i1(inst_doa_i27_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_13 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_14  (
    .i0(inst_doa_i28_006),
    .i1(inst_doa_i29_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_14 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_15  (
    .i0(inst_doa_i30_006),
    .i1(inst_doa_i31_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_15 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_16  (
    .i0(inst_doa_i32_006),
    .i1(inst_doa_i33_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_16 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_17  (
    .i0(inst_doa_i34_006),
    .i1(inst_doa_i35_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_17 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_18  (
    .i0(inst_doa_i36_006),
    .i1(inst_doa_i37_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_18 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_19  (
    .i0(inst_doa_i38_006),
    .i1(inst_doa_i39_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_19 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_2  (
    .i0(inst_doa_i4_006),
    .i1(inst_doa_i5_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_2 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_20  (
    .i0(inst_doa_i40_006),
    .i1(inst_doa_i41_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_20 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_21  (
    .i0(inst_doa_i42_006),
    .i1(inst_doa_i43_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_21 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_22  (
    .i0(inst_doa_i44_006),
    .i1(inst_doa_i45_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_22 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_23  (
    .i0(inst_doa_i46_006),
    .i1(inst_doa_i47_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_23 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_24  (
    .i0(inst_doa_i48_006),
    .i1(inst_doa_i49_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_24 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_25  (
    .i0(inst_doa_i50_006),
    .i1(inst_doa_i51_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_25 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_26  (
    .i0(inst_doa_i52_006),
    .i1(inst_doa_i53_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_26 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_27  (
    .i0(inst_doa_i54_006),
    .i1(inst_doa_i55_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_27 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_28  (
    .i0(inst_doa_i56_006),
    .i1(inst_doa_i57_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_28 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_29  (
    .i0(inst_doa_i58_006),
    .i1(inst_doa_i59_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_29 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_3  (
    .i0(inst_doa_i6_006),
    .i1(inst_doa_i7_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_3 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_30  (
    .i0(inst_doa_i60_006),
    .i1(inst_doa_i61_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_30 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_31  (
    .i0(inst_doa_i62_006),
    .i1(inst_doa_i63_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_31 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_4  (
    .i0(inst_doa_i8_006),
    .i1(inst_doa_i9_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_4 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_5  (
    .i0(inst_doa_i10_006),
    .i1(inst_doa_i11_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_5 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_6  (
    .i0(inst_doa_i12_006),
    .i1(inst_doa_i13_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_6 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_7  (
    .i0(inst_doa_i14_006),
    .i1(inst_doa_i15_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_7 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_8  (
    .i0(inst_doa_i16_006),
    .i1(inst_doa_i17_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_8 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_9  (
    .i0(inst_doa_i18_006),
    .i1(inst_doa_i19_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_9 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b6/B0_0 ),
    .i1(\inst_doa_mux_b6/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_0 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b6/B0_2 ),
    .i1(\inst_doa_mux_b6/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_1 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_10  (
    .i0(\inst_doa_mux_b6/B0_20 ),
    .i1(\inst_doa_mux_b6/B0_21 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_10 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_11  (
    .i0(\inst_doa_mux_b6/B0_22 ),
    .i1(\inst_doa_mux_b6/B0_23 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_11 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_12  (
    .i0(\inst_doa_mux_b6/B0_24 ),
    .i1(\inst_doa_mux_b6/B0_25 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_12 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_13  (
    .i0(\inst_doa_mux_b6/B0_26 ),
    .i1(\inst_doa_mux_b6/B0_27 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_13 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_14  (
    .i0(\inst_doa_mux_b6/B0_28 ),
    .i1(\inst_doa_mux_b6/B0_29 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_14 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_15  (
    .i0(\inst_doa_mux_b6/B0_30 ),
    .i1(\inst_doa_mux_b6/B0_31 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_15 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_2  (
    .i0(\inst_doa_mux_b6/B0_4 ),
    .i1(\inst_doa_mux_b6/B0_5 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_2 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_3  (
    .i0(\inst_doa_mux_b6/B0_6 ),
    .i1(\inst_doa_mux_b6/B0_7 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_3 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_4  (
    .i0(\inst_doa_mux_b6/B0_8 ),
    .i1(\inst_doa_mux_b6/B0_9 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_4 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_5  (
    .i0(\inst_doa_mux_b6/B0_10 ),
    .i1(\inst_doa_mux_b6/B0_11 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_5 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_6  (
    .i0(\inst_doa_mux_b6/B0_12 ),
    .i1(\inst_doa_mux_b6/B0_13 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_6 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_7  (
    .i0(\inst_doa_mux_b6/B0_14 ),
    .i1(\inst_doa_mux_b6/B0_15 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_7 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_8  (
    .i0(\inst_doa_mux_b6/B0_16 ),
    .i1(\inst_doa_mux_b6/B0_17 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_8 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_9  (
    .i0(\inst_doa_mux_b6/B0_18 ),
    .i1(\inst_doa_mux_b6/B0_19 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_9 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b6/B1_0 ),
    .i1(\inst_doa_mux_b6/B1_1 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b6/B2_0 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_2_1  (
    .i0(\inst_doa_mux_b6/B1_2 ),
    .i1(\inst_doa_mux_b6/B1_3 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b6/B2_1 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_2_2  (
    .i0(\inst_doa_mux_b6/B1_4 ),
    .i1(\inst_doa_mux_b6/B1_5 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b6/B2_2 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_2_3  (
    .i0(\inst_doa_mux_b6/B1_6 ),
    .i1(\inst_doa_mux_b6/B1_7 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b6/B2_3 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_2_4  (
    .i0(\inst_doa_mux_b6/B1_8 ),
    .i1(\inst_doa_mux_b6/B1_9 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b6/B2_4 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_2_5  (
    .i0(\inst_doa_mux_b6/B1_10 ),
    .i1(\inst_doa_mux_b6/B1_11 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b6/B2_5 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_2_6  (
    .i0(\inst_doa_mux_b6/B1_12 ),
    .i1(\inst_doa_mux_b6/B1_13 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b6/B2_6 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_2_7  (
    .i0(\inst_doa_mux_b6/B1_14 ),
    .i1(\inst_doa_mux_b6/B1_15 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b6/B2_7 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_3_0  (
    .i0(\inst_doa_mux_b6/B2_0 ),
    .i1(\inst_doa_mux_b6/B2_1 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b6/B3_0 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_3_1  (
    .i0(\inst_doa_mux_b6/B2_2 ),
    .i1(\inst_doa_mux_b6/B2_3 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b6/B3_1 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_3_2  (
    .i0(\inst_doa_mux_b6/B2_4 ),
    .i1(\inst_doa_mux_b6/B2_5 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b6/B3_2 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_3_3  (
    .i0(\inst_doa_mux_b6/B2_6 ),
    .i1(\inst_doa_mux_b6/B2_7 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b6/B3_3 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_4_0  (
    .i0(\inst_doa_mux_b6/B3_0 ),
    .i1(\inst_doa_mux_b6/B3_1 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b6/B4_0 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_4_1  (
    .i0(\inst_doa_mux_b6/B3_2 ),
    .i1(\inst_doa_mux_b6/B3_3 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b6/B4_1 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_5_0  (
    .i0(\inst_doa_mux_b6/B4_0 ),
    .i1(\inst_doa_mux_b6/B4_1 ),
    .sel(addra_piped[5]),
    .o(doa[6]));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_0  (
    .i0(inst_doa_i0_007),
    .i1(inst_doa_i1_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_0 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_1  (
    .i0(inst_doa_i2_007),
    .i1(inst_doa_i3_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_1 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_10  (
    .i0(inst_doa_i20_007),
    .i1(inst_doa_i21_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_10 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_11  (
    .i0(inst_doa_i22_007),
    .i1(inst_doa_i23_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_11 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_12  (
    .i0(inst_doa_i24_007),
    .i1(inst_doa_i25_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_12 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_13  (
    .i0(inst_doa_i26_007),
    .i1(inst_doa_i27_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_13 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_14  (
    .i0(inst_doa_i28_007),
    .i1(inst_doa_i29_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_14 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_15  (
    .i0(inst_doa_i30_007),
    .i1(inst_doa_i31_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_15 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_16  (
    .i0(inst_doa_i32_007),
    .i1(inst_doa_i33_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_16 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_17  (
    .i0(inst_doa_i34_007),
    .i1(inst_doa_i35_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_17 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_18  (
    .i0(inst_doa_i36_007),
    .i1(inst_doa_i37_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_18 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_19  (
    .i0(inst_doa_i38_007),
    .i1(inst_doa_i39_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_19 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_2  (
    .i0(inst_doa_i4_007),
    .i1(inst_doa_i5_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_2 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_20  (
    .i0(inst_doa_i40_007),
    .i1(inst_doa_i41_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_20 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_21  (
    .i0(inst_doa_i42_007),
    .i1(inst_doa_i43_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_21 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_22  (
    .i0(inst_doa_i44_007),
    .i1(inst_doa_i45_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_22 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_23  (
    .i0(inst_doa_i46_007),
    .i1(inst_doa_i47_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_23 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_24  (
    .i0(inst_doa_i48_007),
    .i1(inst_doa_i49_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_24 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_25  (
    .i0(inst_doa_i50_007),
    .i1(inst_doa_i51_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_25 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_26  (
    .i0(inst_doa_i52_007),
    .i1(inst_doa_i53_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_26 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_27  (
    .i0(inst_doa_i54_007),
    .i1(inst_doa_i55_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_27 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_28  (
    .i0(inst_doa_i56_007),
    .i1(inst_doa_i57_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_28 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_29  (
    .i0(inst_doa_i58_007),
    .i1(inst_doa_i59_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_29 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_3  (
    .i0(inst_doa_i6_007),
    .i1(inst_doa_i7_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_3 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_30  (
    .i0(inst_doa_i60_007),
    .i1(inst_doa_i61_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_30 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_31  (
    .i0(inst_doa_i62_007),
    .i1(inst_doa_i63_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_31 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_4  (
    .i0(inst_doa_i8_007),
    .i1(inst_doa_i9_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_4 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_5  (
    .i0(inst_doa_i10_007),
    .i1(inst_doa_i11_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_5 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_6  (
    .i0(inst_doa_i12_007),
    .i1(inst_doa_i13_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_6 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_7  (
    .i0(inst_doa_i14_007),
    .i1(inst_doa_i15_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_7 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_8  (
    .i0(inst_doa_i16_007),
    .i1(inst_doa_i17_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_8 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_9  (
    .i0(inst_doa_i18_007),
    .i1(inst_doa_i19_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_9 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b7/B0_0 ),
    .i1(\inst_doa_mux_b7/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_0 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b7/B0_2 ),
    .i1(\inst_doa_mux_b7/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_1 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_10  (
    .i0(\inst_doa_mux_b7/B0_20 ),
    .i1(\inst_doa_mux_b7/B0_21 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_10 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_11  (
    .i0(\inst_doa_mux_b7/B0_22 ),
    .i1(\inst_doa_mux_b7/B0_23 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_11 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_12  (
    .i0(\inst_doa_mux_b7/B0_24 ),
    .i1(\inst_doa_mux_b7/B0_25 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_12 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_13  (
    .i0(\inst_doa_mux_b7/B0_26 ),
    .i1(\inst_doa_mux_b7/B0_27 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_13 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_14  (
    .i0(\inst_doa_mux_b7/B0_28 ),
    .i1(\inst_doa_mux_b7/B0_29 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_14 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_15  (
    .i0(\inst_doa_mux_b7/B0_30 ),
    .i1(\inst_doa_mux_b7/B0_31 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_15 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_2  (
    .i0(\inst_doa_mux_b7/B0_4 ),
    .i1(\inst_doa_mux_b7/B0_5 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_2 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_3  (
    .i0(\inst_doa_mux_b7/B0_6 ),
    .i1(\inst_doa_mux_b7/B0_7 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_3 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_4  (
    .i0(\inst_doa_mux_b7/B0_8 ),
    .i1(\inst_doa_mux_b7/B0_9 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_4 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_5  (
    .i0(\inst_doa_mux_b7/B0_10 ),
    .i1(\inst_doa_mux_b7/B0_11 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_5 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_6  (
    .i0(\inst_doa_mux_b7/B0_12 ),
    .i1(\inst_doa_mux_b7/B0_13 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_6 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_7  (
    .i0(\inst_doa_mux_b7/B0_14 ),
    .i1(\inst_doa_mux_b7/B0_15 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_7 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_8  (
    .i0(\inst_doa_mux_b7/B0_16 ),
    .i1(\inst_doa_mux_b7/B0_17 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_8 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_9  (
    .i0(\inst_doa_mux_b7/B0_18 ),
    .i1(\inst_doa_mux_b7/B0_19 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_9 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b7/B1_0 ),
    .i1(\inst_doa_mux_b7/B1_1 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b7/B2_0 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_2_1  (
    .i0(\inst_doa_mux_b7/B1_2 ),
    .i1(\inst_doa_mux_b7/B1_3 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b7/B2_1 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_2_2  (
    .i0(\inst_doa_mux_b7/B1_4 ),
    .i1(\inst_doa_mux_b7/B1_5 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b7/B2_2 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_2_3  (
    .i0(\inst_doa_mux_b7/B1_6 ),
    .i1(\inst_doa_mux_b7/B1_7 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b7/B2_3 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_2_4  (
    .i0(\inst_doa_mux_b7/B1_8 ),
    .i1(\inst_doa_mux_b7/B1_9 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b7/B2_4 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_2_5  (
    .i0(\inst_doa_mux_b7/B1_10 ),
    .i1(\inst_doa_mux_b7/B1_11 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b7/B2_5 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_2_6  (
    .i0(\inst_doa_mux_b7/B1_12 ),
    .i1(\inst_doa_mux_b7/B1_13 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b7/B2_6 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_2_7  (
    .i0(\inst_doa_mux_b7/B1_14 ),
    .i1(\inst_doa_mux_b7/B1_15 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b7/B2_7 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_3_0  (
    .i0(\inst_doa_mux_b7/B2_0 ),
    .i1(\inst_doa_mux_b7/B2_1 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b7/B3_0 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_3_1  (
    .i0(\inst_doa_mux_b7/B2_2 ),
    .i1(\inst_doa_mux_b7/B2_3 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b7/B3_1 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_3_2  (
    .i0(\inst_doa_mux_b7/B2_4 ),
    .i1(\inst_doa_mux_b7/B2_5 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b7/B3_2 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_3_3  (
    .i0(\inst_doa_mux_b7/B2_6 ),
    .i1(\inst_doa_mux_b7/B2_7 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b7/B3_3 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_4_0  (
    .i0(\inst_doa_mux_b7/B3_0 ),
    .i1(\inst_doa_mux_b7/B3_1 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b7/B4_0 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_4_1  (
    .i0(\inst_doa_mux_b7/B3_2 ),
    .i1(\inst_doa_mux_b7/B3_3 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b7/B4_1 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_5_0  (
    .i0(\inst_doa_mux_b7/B4_0 ),
    .i1(\inst_doa_mux_b7/B4_1 ),
    .sel(addra_piped[5]),
    .o(doa[7]));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_0  (
    .i0(inst_doa_i0_008),
    .i1(inst_doa_i1_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_0 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_1  (
    .i0(inst_doa_i2_008),
    .i1(inst_doa_i3_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_1 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_10  (
    .i0(inst_doa_i20_008),
    .i1(inst_doa_i21_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_10 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_11  (
    .i0(inst_doa_i22_008),
    .i1(inst_doa_i23_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_11 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_12  (
    .i0(inst_doa_i24_008),
    .i1(inst_doa_i25_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_12 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_13  (
    .i0(inst_doa_i26_008),
    .i1(inst_doa_i27_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_13 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_14  (
    .i0(inst_doa_i28_008),
    .i1(inst_doa_i29_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_14 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_15  (
    .i0(inst_doa_i30_008),
    .i1(inst_doa_i31_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_15 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_16  (
    .i0(inst_doa_i32_008),
    .i1(inst_doa_i33_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_16 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_17  (
    .i0(inst_doa_i34_008),
    .i1(inst_doa_i35_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_17 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_18  (
    .i0(inst_doa_i36_008),
    .i1(inst_doa_i37_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_18 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_19  (
    .i0(inst_doa_i38_008),
    .i1(inst_doa_i39_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_19 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_2  (
    .i0(inst_doa_i4_008),
    .i1(inst_doa_i5_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_2 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_20  (
    .i0(inst_doa_i40_008),
    .i1(inst_doa_i41_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_20 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_21  (
    .i0(inst_doa_i42_008),
    .i1(inst_doa_i43_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_21 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_22  (
    .i0(inst_doa_i44_008),
    .i1(inst_doa_i45_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_22 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_23  (
    .i0(inst_doa_i46_008),
    .i1(inst_doa_i47_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_23 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_24  (
    .i0(inst_doa_i48_008),
    .i1(inst_doa_i49_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_24 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_25  (
    .i0(inst_doa_i50_008),
    .i1(inst_doa_i51_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_25 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_26  (
    .i0(inst_doa_i52_008),
    .i1(inst_doa_i53_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_26 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_27  (
    .i0(inst_doa_i54_008),
    .i1(inst_doa_i55_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_27 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_28  (
    .i0(inst_doa_i56_008),
    .i1(inst_doa_i57_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_28 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_29  (
    .i0(inst_doa_i58_008),
    .i1(inst_doa_i59_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_29 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_3  (
    .i0(inst_doa_i6_008),
    .i1(inst_doa_i7_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_3 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_30  (
    .i0(inst_doa_i60_008),
    .i1(inst_doa_i61_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_30 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_31  (
    .i0(inst_doa_i62_008),
    .i1(inst_doa_i63_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_31 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_4  (
    .i0(inst_doa_i8_008),
    .i1(inst_doa_i9_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_4 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_5  (
    .i0(inst_doa_i10_008),
    .i1(inst_doa_i11_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_5 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_6  (
    .i0(inst_doa_i12_008),
    .i1(inst_doa_i13_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_6 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_7  (
    .i0(inst_doa_i14_008),
    .i1(inst_doa_i15_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_7 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_8  (
    .i0(inst_doa_i16_008),
    .i1(inst_doa_i17_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_8 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_9  (
    .i0(inst_doa_i18_008),
    .i1(inst_doa_i19_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_9 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b8/B0_0 ),
    .i1(\inst_doa_mux_b8/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_0 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b8/B0_2 ),
    .i1(\inst_doa_mux_b8/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_1 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_10  (
    .i0(\inst_doa_mux_b8/B0_20 ),
    .i1(\inst_doa_mux_b8/B0_21 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_10 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_11  (
    .i0(\inst_doa_mux_b8/B0_22 ),
    .i1(\inst_doa_mux_b8/B0_23 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_11 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_12  (
    .i0(\inst_doa_mux_b8/B0_24 ),
    .i1(\inst_doa_mux_b8/B0_25 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_12 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_13  (
    .i0(\inst_doa_mux_b8/B0_26 ),
    .i1(\inst_doa_mux_b8/B0_27 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_13 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_14  (
    .i0(\inst_doa_mux_b8/B0_28 ),
    .i1(\inst_doa_mux_b8/B0_29 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_14 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_15  (
    .i0(\inst_doa_mux_b8/B0_30 ),
    .i1(\inst_doa_mux_b8/B0_31 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_15 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_2  (
    .i0(\inst_doa_mux_b8/B0_4 ),
    .i1(\inst_doa_mux_b8/B0_5 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_2 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_3  (
    .i0(\inst_doa_mux_b8/B0_6 ),
    .i1(\inst_doa_mux_b8/B0_7 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_3 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_4  (
    .i0(\inst_doa_mux_b8/B0_8 ),
    .i1(\inst_doa_mux_b8/B0_9 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_4 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_5  (
    .i0(\inst_doa_mux_b8/B0_10 ),
    .i1(\inst_doa_mux_b8/B0_11 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_5 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_6  (
    .i0(\inst_doa_mux_b8/B0_12 ),
    .i1(\inst_doa_mux_b8/B0_13 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_6 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_7  (
    .i0(\inst_doa_mux_b8/B0_14 ),
    .i1(\inst_doa_mux_b8/B0_15 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_7 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_8  (
    .i0(\inst_doa_mux_b8/B0_16 ),
    .i1(\inst_doa_mux_b8/B0_17 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_8 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_9  (
    .i0(\inst_doa_mux_b8/B0_18 ),
    .i1(\inst_doa_mux_b8/B0_19 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_9 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b8/B1_0 ),
    .i1(\inst_doa_mux_b8/B1_1 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b8/B2_0 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_2_1  (
    .i0(\inst_doa_mux_b8/B1_2 ),
    .i1(\inst_doa_mux_b8/B1_3 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b8/B2_1 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_2_2  (
    .i0(\inst_doa_mux_b8/B1_4 ),
    .i1(\inst_doa_mux_b8/B1_5 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b8/B2_2 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_2_3  (
    .i0(\inst_doa_mux_b8/B1_6 ),
    .i1(\inst_doa_mux_b8/B1_7 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b8/B2_3 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_2_4  (
    .i0(\inst_doa_mux_b8/B1_8 ),
    .i1(\inst_doa_mux_b8/B1_9 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b8/B2_4 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_2_5  (
    .i0(\inst_doa_mux_b8/B1_10 ),
    .i1(\inst_doa_mux_b8/B1_11 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b8/B2_5 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_2_6  (
    .i0(\inst_doa_mux_b8/B1_12 ),
    .i1(\inst_doa_mux_b8/B1_13 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b8/B2_6 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_2_7  (
    .i0(\inst_doa_mux_b8/B1_14 ),
    .i1(\inst_doa_mux_b8/B1_15 ),
    .sel(addra_piped[2]),
    .o(\inst_doa_mux_b8/B2_7 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_3_0  (
    .i0(\inst_doa_mux_b8/B2_0 ),
    .i1(\inst_doa_mux_b8/B2_1 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b8/B3_0 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_3_1  (
    .i0(\inst_doa_mux_b8/B2_2 ),
    .i1(\inst_doa_mux_b8/B2_3 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b8/B3_1 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_3_2  (
    .i0(\inst_doa_mux_b8/B2_4 ),
    .i1(\inst_doa_mux_b8/B2_5 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b8/B3_2 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_3_3  (
    .i0(\inst_doa_mux_b8/B2_6 ),
    .i1(\inst_doa_mux_b8/B2_7 ),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b8/B3_3 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_4_0  (
    .i0(\inst_doa_mux_b8/B3_0 ),
    .i1(\inst_doa_mux_b8/B3_1 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b8/B4_0 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_4_1  (
    .i0(\inst_doa_mux_b8/B3_2 ),
    .i1(\inst_doa_mux_b8/B3_3 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b8/B4_1 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_5_0  (
    .i0(\inst_doa_mux_b8/B4_0 ),
    .i1(\inst_doa_mux_b8/B4_1 ),
    .sel(addra_piped[5]),
    .o(doa[8]));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_3_0  (
    .i0(inst_doa_i0_009),
    .i1(inst_doa_i8_009),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b9/B3_0 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_3_1  (
    .i0(inst_doa_i16_009),
    .i1(inst_doa_i24_009),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b9/B3_1 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_3_2  (
    .i0(inst_doa_i32_009),
    .i1(inst_doa_i40_009),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b9/B3_2 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_3_3  (
    .i0(inst_doa_i48_009),
    .i1(inst_doa_i56_009),
    .sel(addra_piped[3]),
    .o(\inst_doa_mux_b9/B3_3 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_4_0  (
    .i0(\inst_doa_mux_b9/B3_0 ),
    .i1(\inst_doa_mux_b9/B3_1 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b9/B4_0 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_4_1  (
    .i0(\inst_doa_mux_b9/B3_2 ),
    .i1(\inst_doa_mux_b9/B3_3 ),
    .sel(addra_piped[4]),
    .o(\inst_doa_mux_b9/B4_1 ));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_5_0  (
    .i0(\inst_doa_mux_b9/B4_0 ),
    .i1(\inst_doa_mux_b9/B4_1 ),
    .sel(addra_piped[5]),
    .o(doa[9]));

endmodule 

module AL_DFF_X
  (
  ar,
  as,
  clk,
  d,
  en,
  sr,
  ss,
  q
  );

  input ar;
  input as;
  input clk;
  input d;
  input en;
  input sr;
  input ss;
  output q;

  wire enout;
  wire srout;
  wire ssout;

  AL_MUX u_en (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_MUX u_reset (
    .i0(ssout),
    .i1(1'b0),
    .sel(sr),
    .o(srout));
  AL_DFF u_seq (
    .clk(clk),
    .d(srout),
    .reset(ar),
    .set(as),
    .q(q));
  AL_MUX u_set (
    .i0(enout),
    .i1(1'b1),
    .sel(ss),
    .o(ssout));

endmodule 

module AL_MUX
  (
  input i0,
  input i1,
  input sel,
  output o
  );

  wire not_sel, sel_i0, sel_i1;
  not u0 (not_sel, sel);
  and u1 (sel_i1, sel, i1);
  and u2 (sel_i0, not_sel, i0);
  or u3 (o, sel_i1, sel_i0);

endmodule

module AL_DFF
  (
  input reset,
  input set,
  input clk,
  input d,
  output reg q
  );

  parameter INI = 1'b0;

  // synthesis translate_off
  tri0 gsrn = glbl.gsrn;

  always @(gsrn)
  begin
    if(!gsrn)
      assign q = INI;
    else
      deassign q;
  end
  // synthesis translate_on

  always @(posedge reset or posedge set or posedge clk)
  begin
    if (reset)
      q <= 1'b0;
    else if (set)
      q <= 1'b1;
    else
      q <= d;
  end

endmodule

